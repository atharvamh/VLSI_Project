magic
tech scmos
timestamp 1554041646
<< ab >>
rect 29 653 93 725
rect 97 653 129 725
rect 133 653 173 725
rect 177 653 243 725
rect 247 653 303 725
rect 307 653 331 725
rect 491 693 494 730
rect 491 654 494 692
rect 495 689 527 725
rect 495 685 529 689
rect 495 654 527 685
rect 496 653 528 654
rect 533 653 597 725
rect 604 653 676 725
rect 29 581 61 653
rect 65 593 89 653
rect 93 593 133 653
rect 137 593 285 653
rect 494 645 496 653
rect 63 589 285 593
rect 65 581 89 589
rect 93 581 133 589
rect 137 581 285 589
rect 498 581 522 653
rect 530 581 570 653
rect 576 581 608 653
rect 612 581 676 653
rect 29 542 93 581
rect 97 542 129 581
rect 29 538 129 542
rect 29 509 95 538
rect 97 509 129 538
rect 133 509 135 581
rect 137 543 201 581
rect 205 543 259 581
rect 137 539 259 543
rect 137 509 201 539
rect 205 509 259 539
rect 440 509 464 581
rect 466 573 503 581
rect 466 509 503 517
rect 504 509 552 581
rect 556 509 596 581
rect 600 578 624 581
rect 600 510 601 578
rect 602 510 625 578
rect 600 509 624 510
rect 628 509 676 581
rect 29 454 61 509
rect 28 450 61 454
rect 29 436 61 450
rect 65 437 89 509
rect 91 476 133 509
rect 93 439 133 476
rect 93 437 135 439
rect 149 437 213 509
rect 217 439 257 509
rect 217 437 259 439
rect 440 437 504 509
rect 508 437 548 509
rect 552 437 608 509
rect 612 437 676 509
rect 30 416 62 436
rect 28 410 62 416
rect 30 366 62 410
rect 65 366 105 437
rect 109 429 164 437
rect 114 373 154 429
rect 107 367 154 373
rect 156 367 164 373
rect 167 367 207 437
rect 211 367 212 437
rect 24 365 105 366
rect 109 365 165 367
rect 169 365 209 367
rect 213 365 237 437
rect 241 365 281 437
rect 285 365 341 437
rect 416 436 440 437
rect 444 436 484 437
rect 415 365 455 436
rect 460 398 484 436
rect 460 365 485 398
rect 488 365 528 437
rect 532 435 572 437
rect 576 435 632 437
rect 530 365 532 435
rect 536 365 576 435
rect 578 368 632 435
rect 636 368 676 437
rect 578 365 681 368
rect 24 362 127 365
rect 29 293 69 362
rect 73 295 127 362
rect 129 295 169 365
rect 173 295 175 365
rect 73 293 129 295
rect 133 293 173 295
rect 177 293 217 365
rect 220 332 245 365
rect 221 294 245 332
rect 250 294 290 365
rect 221 293 261 294
rect 265 293 289 294
rect 364 293 420 365
rect 424 293 464 365
rect 468 293 492 365
rect 496 363 536 365
rect 540 363 596 365
rect 600 364 681 365
rect 493 293 494 363
rect 498 293 538 363
rect 541 357 549 363
rect 551 357 598 363
rect 551 301 591 357
rect 541 293 596 301
rect 600 293 640 364
rect 643 320 675 364
rect 643 314 677 320
rect 643 294 675 314
rect 29 221 93 293
rect 97 221 153 293
rect 157 221 197 293
rect 201 221 265 293
rect 269 221 293 293
rect 446 291 488 293
rect 448 221 488 291
rect 492 221 556 293
rect 570 291 612 293
rect 572 254 612 291
rect 572 221 614 254
rect 616 221 640 293
rect 644 280 676 294
rect 644 276 677 280
rect 644 221 676 276
rect 29 149 77 221
rect 81 220 105 221
rect 80 152 103 220
rect 104 152 105 220
rect 81 149 105 152
rect 109 149 149 221
rect 153 149 201 221
rect 446 191 500 221
rect 504 191 568 221
rect 446 187 568 191
rect 446 149 500 187
rect 504 149 568 187
rect 570 149 572 221
rect 576 192 608 221
rect 610 192 676 221
rect 576 188 676 192
rect 576 149 608 188
rect 612 149 676 188
rect 29 77 93 149
rect 97 77 129 149
rect 135 77 175 149
rect 183 77 207 149
rect 420 141 568 149
rect 572 141 612 149
rect 616 141 640 149
rect 420 137 642 141
rect 209 77 211 85
rect 420 77 568 137
rect 572 77 612 137
rect 616 77 640 137
rect 644 77 676 149
rect 29 5 101 77
rect 108 5 172 77
rect 177 76 209 77
rect 178 45 210 76
rect 176 41 210 45
rect 178 5 210 41
rect 211 38 214 76
rect 211 0 214 37
rect 374 5 398 77
rect 402 5 458 77
rect 462 5 528 77
rect 532 5 572 77
rect 576 5 608 77
rect 612 5 676 77
<< nwell >>
rect 24 653 336 693
rect 24 613 287 653
rect 491 613 681 693
rect 24 504 262 549
rect 24 469 259 504
rect 435 469 681 549
rect 24 360 341 405
rect 411 370 681 405
rect 24 325 294 360
rect 359 325 681 370
rect 24 216 298 261
rect 446 226 681 261
rect 24 181 206 216
rect 443 181 681 226
rect 24 37 214 117
rect 418 77 681 117
rect 369 37 681 77
<< pwell >>
rect 24 725 330 730
rect 24 693 336 725
rect 491 693 681 730
rect 24 581 287 613
rect 491 586 681 613
rect 24 576 286 581
rect 24 549 262 576
rect 435 549 681 586
rect 24 442 259 469
rect 435 442 681 469
rect 24 405 341 442
rect 411 405 681 442
rect 24 298 294 325
rect 24 261 298 298
rect 359 288 681 325
rect 446 261 681 288
rect 24 154 206 181
rect 443 154 681 181
rect 24 117 214 154
rect 419 149 681 154
rect 418 117 681 149
rect 24 0 214 37
rect 369 5 681 37
rect 375 0 681 5
<< poly >>
rect 41 721 66 723
rect 41 713 43 721
rect 54 713 56 717
rect 64 713 66 721
rect 74 716 76 721
rect 81 716 83 721
rect 38 711 43 713
rect 38 708 40 711
rect 107 713 109 718
rect 118 710 120 714
rect 142 710 144 714
rect 155 712 157 717
rect 162 712 164 717
rect 189 721 214 723
rect 189 713 191 721
rect 202 713 204 717
rect 212 713 214 721
rect 222 716 224 721
rect 229 716 231 721
rect 262 719 264 723
rect 269 719 271 723
rect 276 719 278 723
rect 283 719 285 723
rect 54 701 56 704
rect 47 699 56 701
rect 64 700 66 704
rect 74 701 76 704
rect 38 691 40 699
rect 47 697 49 699
rect 51 697 56 699
rect 47 695 56 697
rect 72 699 76 701
rect 72 696 74 699
rect 54 691 56 695
rect 68 694 74 696
rect 81 695 83 704
rect 107 696 109 705
rect 118 699 120 702
rect 186 711 191 713
rect 186 708 188 711
rect 116 697 122 699
rect 68 692 70 694
rect 72 692 74 694
rect 35 689 48 691
rect 54 689 64 691
rect 68 690 74 692
rect 35 688 37 689
rect 31 686 37 688
rect 46 686 48 689
rect 62 686 64 689
rect 72 686 74 690
rect 78 693 84 695
rect 78 691 80 693
rect 82 691 84 693
rect 78 689 84 691
rect 106 694 112 696
rect 106 692 108 694
rect 110 692 112 694
rect 106 690 112 692
rect 116 695 118 697
rect 120 695 122 697
rect 116 693 122 695
rect 142 696 144 701
rect 155 696 157 701
rect 142 694 148 696
rect 82 686 84 689
rect 109 687 111 690
rect 116 687 118 693
rect 142 692 144 694
rect 146 692 148 694
rect 142 690 148 692
rect 152 694 158 696
rect 152 692 154 694
rect 156 692 158 694
rect 152 690 158 692
rect 31 684 33 686
rect 35 684 37 686
rect 31 682 37 684
rect 62 664 64 668
rect 72 664 74 668
rect 46 655 48 659
rect 142 686 144 690
rect 152 679 154 690
rect 162 688 164 701
rect 202 701 204 704
rect 195 699 204 701
rect 212 700 214 704
rect 222 701 224 704
rect 186 691 188 699
rect 195 697 197 699
rect 199 697 204 699
rect 195 695 204 697
rect 220 699 224 701
rect 220 696 222 699
rect 202 691 204 695
rect 216 694 222 696
rect 229 695 231 704
rect 545 721 570 723
rect 316 708 318 713
rect 505 709 507 714
rect 515 709 517 714
rect 545 713 547 721
rect 558 713 560 717
rect 568 713 570 721
rect 578 716 580 721
rect 585 716 587 721
rect 653 719 655 723
rect 663 719 665 723
rect 542 711 547 713
rect 542 708 544 711
rect 613 708 615 713
rect 558 701 560 704
rect 551 699 560 701
rect 568 700 570 704
rect 578 701 580 704
rect 262 696 264 699
rect 216 692 218 694
rect 220 692 222 694
rect 183 689 196 691
rect 202 689 212 691
rect 216 690 222 692
rect 183 688 185 689
rect 162 686 168 688
rect 162 684 164 686
rect 166 684 168 686
rect 162 682 168 684
rect 179 686 185 688
rect 194 686 196 689
rect 210 686 212 689
rect 220 686 222 690
rect 226 693 232 695
rect 226 691 228 693
rect 230 691 232 693
rect 226 689 232 691
rect 230 686 232 689
rect 256 694 264 696
rect 256 692 258 694
rect 260 693 264 694
rect 260 692 262 693
rect 256 690 262 692
rect 179 684 181 686
rect 183 684 185 686
rect 179 682 185 684
rect 162 679 164 682
rect 142 664 144 668
rect 152 661 154 666
rect 162 661 164 666
rect 82 655 84 659
rect 109 655 111 659
rect 116 655 118 659
rect 210 664 212 668
rect 220 664 222 668
rect 194 655 196 659
rect 256 680 258 690
rect 269 689 271 699
rect 276 689 278 699
rect 283 696 285 699
rect 316 696 318 699
rect 283 694 294 696
rect 286 692 290 694
rect 292 692 294 694
rect 286 690 294 692
rect 316 694 322 696
rect 316 692 318 694
rect 320 692 322 694
rect 316 690 322 692
rect 505 691 507 699
rect 515 695 517 699
rect 515 693 525 695
rect 515 691 521 693
rect 523 691 525 693
rect 542 691 544 699
rect 551 697 553 699
rect 555 697 560 699
rect 551 695 560 697
rect 576 699 580 701
rect 576 696 578 699
rect 558 691 560 695
rect 572 694 578 696
rect 585 695 587 704
rect 637 702 643 704
rect 637 700 639 702
rect 641 700 643 702
rect 613 696 615 699
rect 637 698 643 700
rect 572 692 574 694
rect 576 692 578 694
rect 266 687 272 689
rect 266 685 268 687
rect 270 685 272 687
rect 266 683 272 685
rect 276 687 282 689
rect 276 685 278 687
rect 280 685 282 687
rect 276 683 282 685
rect 266 680 268 683
rect 276 680 278 683
rect 286 680 288 690
rect 316 687 318 690
rect 505 689 525 691
rect 539 689 552 691
rect 558 689 568 691
rect 572 690 578 692
rect 505 684 507 689
rect 515 684 517 689
rect 539 688 541 689
rect 535 686 541 688
rect 550 686 552 689
rect 566 686 568 689
rect 576 686 578 690
rect 582 693 588 695
rect 582 691 584 693
rect 586 691 588 693
rect 582 689 588 691
rect 586 686 588 689
rect 613 694 619 696
rect 613 692 615 694
rect 617 692 619 694
rect 613 690 619 692
rect 613 687 615 690
rect 535 684 537 686
rect 539 684 541 686
rect 316 664 318 669
rect 230 655 232 659
rect 256 658 258 663
rect 266 658 268 663
rect 276 658 278 663
rect 286 658 288 663
rect 535 682 541 684
rect 515 664 517 668
rect 505 656 507 660
rect 566 664 568 668
rect 576 664 578 668
rect 550 655 552 659
rect 641 686 643 698
rect 653 696 655 704
rect 663 701 665 704
rect 648 694 655 696
rect 659 699 665 701
rect 659 697 661 699
rect 663 698 665 699
rect 663 697 667 698
rect 659 695 667 697
rect 648 692 650 694
rect 652 692 655 694
rect 648 691 655 692
rect 648 689 660 691
rect 648 686 650 689
rect 658 686 660 689
rect 665 686 667 695
rect 613 664 615 669
rect 586 655 588 659
rect 641 655 643 659
rect 648 655 650 659
rect 658 655 660 659
rect 665 655 667 659
rect 38 647 40 651
rect 48 647 50 651
rect 74 637 76 642
rect 102 638 104 642
rect 112 640 114 645
rect 122 640 124 645
rect 38 616 40 623
rect 48 620 50 623
rect 48 618 59 620
rect 146 639 148 644
rect 156 639 158 644
rect 166 639 168 644
rect 218 645 220 650
rect 225 645 227 650
rect 232 645 234 650
rect 239 645 241 650
rect 48 616 55 618
rect 57 616 59 618
rect 38 614 44 616
rect 38 612 40 614
rect 42 612 44 614
rect 38 610 44 612
rect 48 614 59 616
rect 74 616 76 619
rect 102 616 104 620
rect 112 616 114 627
rect 122 624 124 627
rect 122 622 128 624
rect 122 620 124 622
rect 126 620 128 622
rect 178 638 180 643
rect 122 618 128 620
rect 74 614 80 616
rect 41 607 43 610
rect 48 607 50 614
rect 74 612 76 614
rect 78 612 80 614
rect 74 610 80 612
rect 102 614 108 616
rect 102 612 104 614
rect 106 612 108 614
rect 102 610 108 612
rect 112 614 118 616
rect 112 612 114 614
rect 116 612 118 614
rect 112 610 118 612
rect 74 607 76 610
rect 102 605 104 610
rect 115 605 117 610
rect 122 605 124 618
rect 146 616 148 621
rect 156 616 158 626
rect 166 623 168 626
rect 166 621 172 623
rect 166 619 168 621
rect 170 619 172 621
rect 166 617 172 619
rect 146 614 152 616
rect 146 612 148 614
rect 150 612 152 614
rect 146 610 152 612
rect 156 614 162 616
rect 156 612 158 614
rect 160 612 162 614
rect 156 610 162 612
rect 146 606 148 610
rect 159 606 161 610
rect 166 606 168 617
rect 178 616 180 625
rect 587 647 589 651
rect 597 647 599 651
rect 621 647 623 651
rect 249 638 251 642
rect 256 638 258 642
rect 263 638 265 642
rect 270 638 272 642
rect 511 637 513 642
rect 539 638 541 642
rect 549 640 551 645
rect 559 640 561 645
rect 218 617 220 620
rect 178 614 184 616
rect 178 612 180 614
rect 182 612 184 614
rect 173 610 184 612
rect 207 615 220 617
rect 207 613 209 615
rect 211 613 216 615
rect 207 611 216 613
rect 173 606 175 610
rect 74 593 76 598
rect 102 592 104 596
rect 41 583 43 587
rect 48 583 50 587
rect 115 589 117 594
rect 122 589 124 594
rect 146 592 148 597
rect 214 599 216 611
rect 225 610 227 620
rect 232 617 234 620
rect 239 617 241 620
rect 249 617 251 620
rect 232 614 235 617
rect 239 615 251 617
rect 222 608 228 610
rect 222 606 224 608
rect 226 606 228 608
rect 222 604 228 606
rect 233 608 235 614
rect 233 606 239 608
rect 233 604 235 606
rect 237 604 239 606
rect 224 599 226 604
rect 233 602 239 604
rect 236 599 238 602
rect 246 599 248 615
rect 256 608 258 620
rect 263 611 265 620
rect 270 617 272 620
rect 270 615 278 617
rect 511 616 513 619
rect 272 613 274 615
rect 276 613 278 615
rect 272 611 278 613
rect 507 614 513 616
rect 507 612 509 614
rect 511 612 513 614
rect 252 606 258 608
rect 252 604 254 606
rect 256 604 258 606
rect 262 609 268 611
rect 507 610 513 612
rect 262 607 264 609
rect 266 607 268 609
rect 511 607 513 610
rect 539 616 541 620
rect 549 616 551 627
rect 559 624 561 627
rect 559 622 565 624
rect 559 620 561 622
rect 563 620 565 622
rect 587 620 589 623
rect 559 618 565 620
rect 578 618 589 620
rect 539 614 545 616
rect 539 612 541 614
rect 543 612 545 614
rect 539 610 545 612
rect 549 614 555 616
rect 549 612 551 614
rect 553 612 555 614
rect 549 610 555 612
rect 262 605 268 607
rect 252 602 258 604
rect 262 598 268 600
rect 262 596 264 598
rect 266 596 268 598
rect 262 594 268 596
rect 159 588 161 593
rect 166 588 168 593
rect 173 588 175 593
rect 214 588 216 593
rect 224 588 226 593
rect 236 588 238 593
rect 246 590 248 593
rect 262 590 264 594
rect 246 588 264 590
rect 539 605 541 610
rect 552 605 554 610
rect 559 605 561 618
rect 578 616 580 618
rect 582 616 589 618
rect 597 616 599 623
rect 657 647 659 651
rect 631 638 633 642
rect 641 638 643 642
rect 668 622 674 624
rect 668 620 670 622
rect 672 620 674 622
rect 578 614 589 616
rect 587 607 589 614
rect 593 614 599 616
rect 593 612 595 614
rect 597 612 599 614
rect 593 610 599 612
rect 621 617 623 620
rect 621 615 627 617
rect 621 613 623 615
rect 625 613 627 615
rect 621 611 627 613
rect 631 616 633 620
rect 641 617 643 620
rect 657 617 659 620
rect 668 618 674 620
rect 668 617 670 618
rect 631 614 637 616
rect 641 615 651 617
rect 657 615 670 617
rect 631 612 633 614
rect 635 612 637 614
rect 594 607 596 610
rect 511 593 513 598
rect 539 592 541 596
rect 552 589 554 594
rect 559 589 561 594
rect 622 602 624 611
rect 631 610 637 612
rect 649 611 651 615
rect 631 607 633 610
rect 629 605 633 607
rect 649 609 658 611
rect 649 607 654 609
rect 656 607 658 609
rect 665 607 667 615
rect 629 602 631 605
rect 639 602 641 606
rect 649 605 658 607
rect 649 602 651 605
rect 665 595 667 598
rect 662 593 667 595
rect 587 583 589 587
rect 594 583 596 587
rect 622 585 624 590
rect 629 585 631 590
rect 639 585 641 593
rect 649 589 651 593
rect 662 585 664 593
rect 639 583 664 585
rect 41 577 66 579
rect 41 569 43 577
rect 54 569 56 573
rect 64 569 66 577
rect 74 572 76 577
rect 81 572 83 577
rect 109 575 111 579
rect 116 575 118 579
rect 38 567 43 569
rect 38 564 40 567
rect 54 557 56 560
rect 47 555 56 557
rect 64 556 66 560
rect 74 557 76 560
rect 38 547 40 555
rect 47 553 49 555
rect 51 553 56 555
rect 47 551 56 553
rect 72 555 76 557
rect 72 552 74 555
rect 54 547 56 551
rect 68 550 74 552
rect 81 551 83 560
rect 168 573 170 578
rect 178 573 180 578
rect 190 573 192 578
rect 223 569 225 574
rect 230 569 232 574
rect 237 569 239 574
rect 529 575 531 579
rect 539 575 541 579
rect 168 560 170 563
rect 178 560 180 563
rect 190 560 192 563
rect 164 558 170 560
rect 153 556 159 558
rect 109 552 111 555
rect 68 548 70 550
rect 72 548 74 550
rect 35 545 48 547
rect 54 545 64 547
rect 68 546 74 548
rect 35 544 37 545
rect 31 542 37 544
rect 46 542 48 545
rect 62 542 64 545
rect 72 542 74 546
rect 78 549 84 551
rect 78 547 80 549
rect 82 547 84 549
rect 78 545 84 547
rect 82 542 84 545
rect 106 550 112 552
rect 106 548 108 550
rect 110 548 112 550
rect 106 546 112 548
rect 116 548 118 555
rect 153 554 155 556
rect 157 554 159 556
rect 153 552 159 554
rect 143 550 149 552
rect 143 548 145 550
rect 147 548 149 550
rect 116 546 127 548
rect 143 546 152 548
rect 31 540 33 542
rect 35 540 37 542
rect 31 538 37 540
rect 62 520 64 524
rect 72 520 74 524
rect 46 511 48 515
rect 106 539 108 546
rect 116 544 123 546
rect 125 544 127 546
rect 116 542 127 544
rect 150 543 152 546
rect 157 543 159 552
rect 164 556 166 558
rect 168 556 170 558
rect 164 554 170 556
rect 176 558 182 560
rect 176 556 178 558
rect 180 556 182 558
rect 176 554 182 556
rect 186 558 192 560
rect 186 556 188 558
rect 190 556 192 558
rect 250 565 252 570
rect 449 564 451 569
rect 186 554 192 556
rect 164 548 166 554
rect 180 549 182 554
rect 164 546 176 548
rect 180 546 183 549
rect 164 543 166 546
rect 174 543 176 546
rect 181 543 183 546
rect 188 543 190 554
rect 223 552 225 556
rect 214 550 225 552
rect 214 548 216 550
rect 218 548 220 550
rect 214 546 220 548
rect 116 539 118 542
rect 218 537 220 546
rect 230 545 232 556
rect 237 552 239 556
rect 250 552 252 556
rect 565 568 567 573
rect 572 568 574 573
rect 653 575 655 579
rect 663 575 665 579
rect 513 558 519 560
rect 513 556 515 558
rect 517 556 519 558
rect 236 550 242 552
rect 236 548 238 550
rect 240 548 242 550
rect 236 546 242 548
rect 246 550 252 552
rect 246 548 248 550
rect 250 548 252 550
rect 246 546 252 548
rect 226 543 232 545
rect 226 541 228 543
rect 230 541 232 543
rect 226 539 232 541
rect 230 536 232 539
rect 240 536 242 546
rect 250 541 252 546
rect 449 552 451 555
rect 513 554 519 556
rect 449 550 455 552
rect 449 548 451 550
rect 453 548 455 550
rect 449 546 455 548
rect 449 543 451 546
rect 218 519 220 524
rect 517 542 519 554
rect 529 552 531 560
rect 539 557 541 560
rect 585 566 587 570
rect 611 564 613 569
rect 524 550 531 552
rect 535 555 541 557
rect 535 553 537 555
rect 539 554 541 555
rect 539 553 543 554
rect 535 551 543 553
rect 524 548 526 550
rect 528 548 531 550
rect 524 547 531 548
rect 524 545 536 547
rect 524 542 526 545
rect 534 542 536 545
rect 541 542 543 551
rect 565 544 567 557
rect 572 552 574 557
rect 585 552 587 557
rect 637 558 643 560
rect 637 556 639 558
rect 641 556 643 558
rect 571 550 577 552
rect 571 548 573 550
rect 575 548 577 550
rect 571 546 577 548
rect 581 550 587 552
rect 581 548 583 550
rect 585 548 587 550
rect 581 546 587 548
rect 561 542 567 544
rect 82 511 84 515
rect 106 511 108 515
rect 116 511 118 515
rect 150 511 152 515
rect 157 511 159 515
rect 164 511 166 515
rect 174 511 176 515
rect 181 511 183 515
rect 188 511 190 515
rect 230 518 232 523
rect 240 518 242 523
rect 250 518 252 523
rect 449 520 451 525
rect 561 540 563 542
rect 565 540 567 542
rect 561 538 567 540
rect 565 535 567 538
rect 575 535 577 546
rect 585 542 587 546
rect 611 552 613 555
rect 637 554 643 556
rect 611 550 617 552
rect 611 548 613 550
rect 615 548 617 550
rect 611 546 617 548
rect 611 543 613 546
rect 641 542 643 554
rect 653 552 655 560
rect 663 557 665 560
rect 648 550 655 552
rect 659 555 665 557
rect 659 553 661 555
rect 663 554 665 555
rect 663 553 667 554
rect 659 551 667 553
rect 648 548 650 550
rect 652 548 655 550
rect 648 547 655 548
rect 648 545 660 547
rect 648 542 650 545
rect 658 542 660 545
rect 665 542 667 551
rect 565 517 567 522
rect 575 517 577 522
rect 585 520 587 524
rect 611 520 613 525
rect 517 511 519 515
rect 524 511 526 515
rect 534 511 536 515
rect 541 511 543 515
rect 641 511 643 515
rect 648 511 650 515
rect 658 511 660 515
rect 665 511 667 515
rect 41 503 43 507
rect 48 503 50 507
rect 158 503 160 507
rect 74 493 76 498
rect 102 494 104 498
rect 112 496 114 501
rect 122 496 124 501
rect 41 472 43 475
rect 38 470 44 472
rect 38 468 40 470
rect 42 468 44 470
rect 38 466 44 468
rect 48 469 50 475
rect 74 472 76 475
rect 102 472 104 476
rect 112 472 114 483
rect 122 480 124 483
rect 122 478 128 480
rect 122 476 124 478
rect 126 476 128 478
rect 194 503 196 507
rect 168 494 170 498
rect 178 494 180 498
rect 449 503 451 507
rect 226 496 228 501
rect 236 496 238 501
rect 246 494 248 498
rect 226 480 228 483
rect 205 478 211 480
rect 205 476 207 478
rect 209 476 211 478
rect 122 474 128 476
rect 74 470 80 472
rect 48 467 54 469
rect 39 457 41 466
rect 48 465 50 467
rect 52 465 54 467
rect 48 463 54 465
rect 74 468 76 470
rect 78 468 80 470
rect 74 466 80 468
rect 102 470 108 472
rect 102 468 104 470
rect 106 468 108 470
rect 102 466 108 468
rect 112 470 118 472
rect 112 468 114 470
rect 116 468 118 470
rect 112 466 118 468
rect 74 463 76 466
rect 50 460 52 463
rect 102 461 104 466
rect 115 461 117 466
rect 122 461 124 474
rect 158 473 160 476
rect 158 471 164 473
rect 158 469 160 471
rect 162 469 164 471
rect 158 467 164 469
rect 168 472 170 476
rect 178 473 180 476
rect 194 473 196 476
rect 205 474 211 476
rect 222 478 228 480
rect 222 476 224 478
rect 226 476 228 478
rect 222 474 228 476
rect 205 473 207 474
rect 168 470 174 472
rect 178 471 188 473
rect 194 471 207 473
rect 168 468 170 470
rect 172 468 174 470
rect 39 444 41 449
rect 50 448 52 452
rect 74 449 76 454
rect 102 448 104 452
rect 159 458 161 467
rect 168 466 174 468
rect 186 467 188 471
rect 168 463 170 466
rect 166 461 170 463
rect 186 465 195 467
rect 186 463 191 465
rect 193 463 195 465
rect 202 463 204 471
rect 166 458 168 461
rect 176 458 178 462
rect 186 461 195 463
rect 186 458 188 461
rect 115 445 117 450
rect 122 445 124 450
rect 226 461 228 474
rect 236 472 238 483
rect 485 503 487 507
rect 459 494 461 498
rect 469 494 471 498
rect 621 503 623 507
rect 517 494 519 498
rect 527 496 529 501
rect 537 496 539 501
rect 496 478 502 480
rect 496 476 498 478
rect 500 476 502 478
rect 562 494 564 498
rect 572 494 574 499
rect 582 494 584 499
rect 592 494 594 499
rect 246 472 248 476
rect 232 470 238 472
rect 232 468 234 470
rect 236 468 238 470
rect 232 466 238 468
rect 242 470 248 472
rect 242 468 244 470
rect 246 468 248 470
rect 242 466 248 468
rect 449 473 451 476
rect 449 471 455 473
rect 449 469 451 471
rect 453 469 455 471
rect 449 467 455 469
rect 459 472 461 476
rect 469 473 471 476
rect 485 473 487 476
rect 496 474 502 476
rect 496 473 498 474
rect 459 470 465 472
rect 469 471 479 473
rect 485 471 498 473
rect 517 472 519 476
rect 527 472 529 483
rect 537 480 539 483
rect 537 478 543 480
rect 537 476 539 478
rect 541 476 543 478
rect 657 503 659 507
rect 631 494 633 498
rect 641 494 643 498
rect 668 478 674 480
rect 668 476 670 478
rect 672 476 674 478
rect 537 474 543 476
rect 459 468 461 470
rect 463 468 465 470
rect 233 461 235 466
rect 246 461 248 466
rect 202 451 204 454
rect 199 449 204 451
rect 450 458 452 467
rect 459 466 465 468
rect 477 467 479 471
rect 459 463 461 466
rect 457 461 461 463
rect 477 465 486 467
rect 477 463 482 465
rect 484 463 486 465
rect 493 463 495 471
rect 517 470 523 472
rect 517 468 519 470
rect 521 468 523 470
rect 517 466 523 468
rect 527 470 533 472
rect 527 468 529 470
rect 531 468 533 470
rect 527 466 533 468
rect 457 458 459 461
rect 467 458 469 462
rect 477 461 486 463
rect 477 458 479 461
rect 159 441 161 446
rect 166 441 168 446
rect 176 441 178 449
rect 186 445 188 449
rect 199 441 201 449
rect 176 439 201 441
rect 226 445 228 450
rect 233 445 235 450
rect 246 448 248 452
rect 517 461 519 466
rect 530 461 532 466
rect 537 461 539 474
rect 562 472 564 476
rect 572 472 574 476
rect 561 470 574 472
rect 561 468 563 470
rect 565 468 574 470
rect 561 466 574 468
rect 561 463 563 466
rect 572 463 574 466
rect 582 472 584 476
rect 592 472 594 476
rect 621 473 623 476
rect 582 470 599 472
rect 582 468 595 470
rect 597 468 599 470
rect 582 466 599 468
rect 621 471 627 473
rect 621 469 623 471
rect 625 469 627 471
rect 621 467 627 469
rect 631 472 633 476
rect 641 473 643 476
rect 657 473 659 476
rect 668 474 674 476
rect 668 473 670 474
rect 631 470 637 472
rect 641 471 651 473
rect 657 471 670 473
rect 631 468 633 470
rect 635 468 637 470
rect 582 463 584 466
rect 592 463 594 466
rect 493 451 495 454
rect 490 449 495 451
rect 450 441 452 446
rect 457 441 459 446
rect 467 441 469 449
rect 477 445 479 449
rect 490 441 492 449
rect 517 448 519 452
rect 467 439 492 441
rect 530 445 532 450
rect 537 445 539 450
rect 561 448 563 452
rect 622 458 624 467
rect 631 466 637 468
rect 649 467 651 471
rect 631 463 633 466
rect 629 461 633 463
rect 649 465 658 467
rect 649 463 654 465
rect 656 463 658 465
rect 665 463 667 471
rect 629 458 631 461
rect 639 458 641 462
rect 649 461 658 463
rect 649 458 651 461
rect 572 439 574 444
rect 582 443 584 448
rect 592 443 594 448
rect 665 451 667 454
rect 662 449 667 451
rect 622 441 624 446
rect 629 441 631 446
rect 639 441 641 449
rect 649 445 651 449
rect 662 441 664 449
rect 639 439 664 441
rect 44 430 46 435
rect 51 430 53 435
rect 74 422 76 426
rect 87 424 89 429
rect 94 424 96 429
rect 44 415 46 418
rect 36 413 46 415
rect 36 411 38 413
rect 40 411 42 413
rect 36 409 42 411
rect 40 394 42 409
rect 51 408 53 418
rect 123 422 125 426
rect 136 424 138 429
rect 143 424 145 429
rect 176 424 178 429
rect 183 424 185 429
rect 196 422 198 426
rect 222 420 224 425
rect 250 422 252 426
rect 263 424 265 429
rect 270 424 272 429
rect 47 406 53 408
rect 47 404 49 406
rect 51 404 53 406
rect 47 402 53 404
rect 74 408 76 413
rect 87 408 89 413
rect 74 406 80 408
rect 74 404 76 406
rect 78 404 80 406
rect 74 402 80 404
rect 84 406 90 408
rect 84 404 86 406
rect 88 404 90 406
rect 84 402 90 404
rect 50 394 52 402
rect 74 398 76 402
rect 84 391 86 402
rect 94 400 96 413
rect 123 408 125 413
rect 136 408 138 413
rect 123 406 129 408
rect 123 404 125 406
rect 127 404 129 406
rect 123 402 129 404
rect 133 406 139 408
rect 133 404 135 406
rect 137 404 139 406
rect 133 402 139 404
rect 94 398 100 400
rect 123 398 125 402
rect 94 396 96 398
rect 98 396 100 398
rect 94 394 100 396
rect 94 391 96 394
rect 40 376 42 380
rect 50 375 52 380
rect 74 376 76 380
rect 133 391 135 402
rect 143 400 145 413
rect 176 400 178 413
rect 183 408 185 413
rect 196 408 198 413
rect 294 421 296 426
rect 307 425 309 430
rect 314 425 316 430
rect 321 425 323 430
rect 182 406 188 408
rect 182 404 184 406
rect 186 404 188 406
rect 182 402 188 404
rect 192 406 198 408
rect 192 404 194 406
rect 196 404 198 406
rect 192 402 198 404
rect 143 398 149 400
rect 143 396 145 398
rect 147 396 149 398
rect 143 394 149 396
rect 172 398 178 400
rect 172 396 174 398
rect 176 396 178 398
rect 172 394 178 396
rect 143 391 145 394
rect 176 391 178 394
rect 186 391 188 402
rect 196 398 198 402
rect 222 408 224 411
rect 250 408 252 413
rect 263 408 265 413
rect 222 406 228 408
rect 222 404 224 406
rect 226 404 228 406
rect 222 402 228 404
rect 250 406 256 408
rect 250 404 252 406
rect 254 404 256 406
rect 250 402 256 404
rect 260 406 266 408
rect 260 404 262 406
rect 264 404 266 406
rect 260 402 266 404
rect 222 399 224 402
rect 84 373 86 378
rect 94 373 96 378
rect 123 376 125 380
rect 250 398 252 402
rect 133 373 135 378
rect 143 373 145 378
rect 176 373 178 378
rect 186 373 188 378
rect 196 376 198 380
rect 222 376 224 381
rect 260 391 262 402
rect 270 400 272 413
rect 424 424 426 429
rect 431 424 433 429
rect 444 422 446 426
rect 469 420 471 425
rect 497 424 499 429
rect 504 424 506 429
rect 294 408 296 412
rect 307 408 309 412
rect 294 406 300 408
rect 294 404 296 406
rect 298 404 300 406
rect 294 402 300 404
rect 304 406 310 408
rect 304 404 306 406
rect 308 404 310 406
rect 304 402 310 404
rect 270 398 276 400
rect 270 396 272 398
rect 274 396 276 398
rect 294 397 296 402
rect 270 394 276 396
rect 270 391 272 394
rect 250 376 252 380
rect 304 392 306 402
rect 314 401 316 412
rect 321 408 323 412
rect 321 406 332 408
rect 326 404 328 406
rect 330 404 332 406
rect 326 402 332 404
rect 314 399 320 401
rect 314 397 316 399
rect 318 397 320 399
rect 314 395 320 397
rect 314 392 316 395
rect 326 393 328 402
rect 424 400 426 413
rect 431 408 433 413
rect 444 408 446 413
rect 517 422 519 426
rect 545 422 547 426
rect 558 424 560 429
rect 565 424 567 429
rect 594 425 596 430
rect 601 425 603 430
rect 608 425 610 430
rect 648 431 650 435
rect 655 431 657 435
rect 662 431 664 435
rect 430 406 436 408
rect 430 404 432 406
rect 434 404 436 406
rect 430 402 436 404
rect 440 406 446 408
rect 440 404 442 406
rect 444 404 446 406
rect 440 402 446 404
rect 420 398 426 400
rect 420 396 422 398
rect 424 396 426 398
rect 420 394 426 396
rect 424 391 426 394
rect 434 391 436 402
rect 444 398 446 402
rect 469 408 471 411
rect 469 406 475 408
rect 469 404 471 406
rect 473 404 475 406
rect 469 402 475 404
rect 469 399 471 402
rect 497 400 499 413
rect 504 408 506 413
rect 517 408 519 413
rect 503 406 509 408
rect 503 404 505 406
rect 507 404 509 406
rect 503 402 509 404
rect 513 406 519 408
rect 513 404 515 406
rect 517 404 519 406
rect 513 402 519 404
rect 260 373 262 378
rect 270 373 272 378
rect 294 374 296 379
rect 304 374 306 379
rect 314 374 316 379
rect 326 375 328 380
rect 493 398 499 400
rect 493 396 495 398
rect 497 396 499 398
rect 493 394 499 396
rect 497 391 499 394
rect 507 391 509 402
rect 517 398 519 402
rect 545 408 547 413
rect 558 408 560 413
rect 545 406 551 408
rect 545 404 547 406
rect 549 404 551 406
rect 545 402 551 404
rect 555 406 561 408
rect 555 404 557 406
rect 559 404 561 406
rect 555 402 561 404
rect 545 398 547 402
rect 424 373 426 378
rect 434 373 436 378
rect 444 376 446 380
rect 469 376 471 381
rect 555 391 557 402
rect 565 400 567 413
rect 621 421 623 426
rect 594 408 596 412
rect 585 406 596 408
rect 585 404 587 406
rect 589 404 591 406
rect 585 402 591 404
rect 565 398 571 400
rect 565 396 567 398
rect 569 396 571 398
rect 565 394 571 396
rect 565 391 567 394
rect 589 393 591 402
rect 601 401 603 412
rect 608 408 610 412
rect 621 408 623 412
rect 648 408 650 411
rect 607 406 613 408
rect 607 404 609 406
rect 611 404 613 406
rect 607 402 613 404
rect 617 406 623 408
rect 617 404 619 406
rect 621 404 623 406
rect 617 402 623 404
rect 641 406 650 408
rect 641 404 643 406
rect 645 404 647 406
rect 641 402 647 404
rect 597 399 603 401
rect 597 397 599 399
rect 601 397 603 399
rect 597 395 603 397
rect 497 373 499 378
rect 507 373 509 378
rect 517 376 519 380
rect 545 376 547 380
rect 601 392 603 395
rect 611 392 613 402
rect 621 397 623 402
rect 555 373 557 378
rect 565 373 567 378
rect 589 375 591 380
rect 645 391 647 402
rect 655 400 657 411
rect 662 408 664 411
rect 661 406 667 408
rect 661 404 663 406
rect 665 404 667 406
rect 661 402 667 404
rect 651 398 657 400
rect 651 396 653 398
rect 655 396 657 398
rect 651 394 657 396
rect 655 391 657 394
rect 665 391 667 402
rect 601 374 603 379
rect 611 374 613 379
rect 621 374 623 379
rect 645 367 647 371
rect 655 367 657 371
rect 665 367 667 371
rect 38 359 40 363
rect 48 359 50 363
rect 58 359 60 363
rect 82 351 84 356
rect 92 351 94 356
rect 102 351 104 356
rect 38 328 40 339
rect 48 336 50 339
rect 48 334 54 336
rect 48 332 50 334
rect 52 332 54 334
rect 48 330 54 332
rect 38 326 44 328
rect 38 324 40 326
rect 42 324 44 326
rect 38 322 44 324
rect 41 319 43 322
rect 48 319 50 330
rect 58 328 60 339
rect 114 350 116 355
rect 138 352 140 357
rect 148 352 150 357
rect 82 328 84 333
rect 92 328 94 338
rect 102 335 104 338
rect 158 350 160 354
rect 186 350 188 354
rect 196 352 198 357
rect 206 352 208 357
rect 102 333 108 335
rect 102 331 104 333
rect 106 331 108 333
rect 102 329 108 331
rect 58 326 64 328
rect 58 324 60 326
rect 62 324 64 326
rect 55 322 64 324
rect 82 326 88 328
rect 82 324 84 326
rect 86 324 88 326
rect 82 322 88 324
rect 92 326 98 328
rect 92 324 94 326
rect 96 324 98 326
rect 92 322 98 324
rect 55 319 57 322
rect 82 318 84 322
rect 95 318 97 322
rect 102 318 104 329
rect 114 328 116 337
rect 138 336 140 339
rect 134 334 140 336
rect 134 332 136 334
rect 138 332 140 334
rect 134 330 140 332
rect 114 326 120 328
rect 114 324 116 326
rect 118 324 120 326
rect 109 322 120 324
rect 109 318 111 322
rect 82 304 84 309
rect 138 317 140 330
rect 148 328 150 339
rect 234 349 236 354
rect 259 350 261 354
rect 269 352 271 357
rect 279 352 281 357
rect 158 328 160 332
rect 144 326 150 328
rect 144 324 146 326
rect 148 324 150 326
rect 144 322 150 324
rect 154 326 160 328
rect 154 324 156 326
rect 158 324 160 326
rect 154 322 160 324
rect 145 317 147 322
rect 158 317 160 322
rect 186 328 188 332
rect 196 328 198 339
rect 206 336 208 339
rect 206 334 212 336
rect 206 332 208 334
rect 210 332 212 334
rect 206 330 212 332
rect 377 350 379 355
rect 389 351 391 356
rect 399 351 401 356
rect 409 351 411 356
rect 433 352 435 357
rect 443 352 445 357
rect 186 326 192 328
rect 186 324 188 326
rect 190 324 192 326
rect 186 322 192 324
rect 196 326 202 328
rect 196 324 198 326
rect 200 324 202 326
rect 196 322 202 324
rect 186 317 188 322
rect 199 317 201 322
rect 206 317 208 330
rect 234 328 236 331
rect 230 326 236 328
rect 230 324 232 326
rect 234 324 236 326
rect 230 322 236 324
rect 234 319 236 322
rect 259 328 261 332
rect 269 328 271 339
rect 279 336 281 339
rect 279 334 285 336
rect 279 332 281 334
rect 283 332 285 334
rect 279 330 285 332
rect 259 326 265 328
rect 259 324 261 326
rect 263 324 265 326
rect 259 322 265 324
rect 269 326 275 328
rect 269 324 271 326
rect 273 324 275 326
rect 269 322 275 324
rect 41 295 43 299
rect 48 295 50 299
rect 55 295 57 299
rect 95 300 97 305
rect 102 300 104 305
rect 109 300 111 305
rect 138 301 140 306
rect 145 301 147 306
rect 158 304 160 308
rect 186 304 188 308
rect 259 317 261 322
rect 272 317 274 322
rect 279 317 281 330
rect 377 328 379 337
rect 389 335 391 338
rect 385 333 391 335
rect 385 331 387 333
rect 389 331 391 333
rect 385 329 391 331
rect 373 326 379 328
rect 373 324 375 326
rect 377 324 379 326
rect 373 322 384 324
rect 382 318 384 322
rect 389 318 391 329
rect 399 328 401 338
rect 453 350 455 354
rect 433 336 435 339
rect 429 334 435 336
rect 409 328 411 333
rect 429 332 431 334
rect 433 332 435 334
rect 429 330 435 332
rect 395 326 401 328
rect 395 324 397 326
rect 399 324 401 326
rect 395 322 401 324
rect 405 326 411 328
rect 405 324 407 326
rect 409 324 411 326
rect 405 322 411 324
rect 396 318 398 322
rect 409 318 411 322
rect 199 301 201 306
rect 206 301 208 306
rect 234 305 236 310
rect 259 304 261 308
rect 272 301 274 306
rect 279 301 281 306
rect 433 317 435 330
rect 443 328 445 339
rect 481 349 483 354
rect 507 350 509 354
rect 517 352 519 357
rect 527 352 529 357
rect 560 352 562 357
rect 570 352 572 357
rect 453 328 455 332
rect 580 350 582 354
rect 609 352 611 357
rect 619 352 621 357
rect 481 328 483 331
rect 439 326 445 328
rect 439 324 441 326
rect 443 324 445 326
rect 439 322 445 324
rect 449 326 455 328
rect 449 324 451 326
rect 453 324 455 326
rect 449 322 455 324
rect 477 326 483 328
rect 477 324 479 326
rect 481 324 483 326
rect 477 322 483 324
rect 440 317 442 322
rect 453 317 455 322
rect 481 319 483 322
rect 507 328 509 332
rect 517 328 519 339
rect 527 336 529 339
rect 560 336 562 339
rect 527 334 533 336
rect 527 332 529 334
rect 531 332 533 334
rect 527 330 533 332
rect 556 334 562 336
rect 556 332 558 334
rect 560 332 562 334
rect 556 330 562 332
rect 507 326 513 328
rect 507 324 509 326
rect 511 324 513 326
rect 507 322 513 324
rect 517 326 523 328
rect 517 324 519 326
rect 521 324 523 326
rect 517 322 523 324
rect 382 300 384 305
rect 389 300 391 305
rect 396 300 398 305
rect 409 304 411 309
rect 507 317 509 322
rect 520 317 522 322
rect 527 317 529 330
rect 560 317 562 330
rect 570 328 572 339
rect 629 350 631 354
rect 653 350 655 355
rect 663 350 665 354
rect 609 336 611 339
rect 605 334 611 336
rect 605 332 607 334
rect 609 332 611 334
rect 580 328 582 332
rect 605 330 611 332
rect 566 326 572 328
rect 566 324 568 326
rect 570 324 572 326
rect 566 322 572 324
rect 576 326 582 328
rect 576 324 578 326
rect 580 324 582 326
rect 576 322 582 324
rect 567 317 569 322
rect 580 317 582 322
rect 609 317 611 330
rect 619 328 621 339
rect 629 328 631 332
rect 653 328 655 336
rect 615 326 621 328
rect 615 324 617 326
rect 619 324 621 326
rect 615 322 621 324
rect 625 326 631 328
rect 625 324 627 326
rect 629 324 631 326
rect 625 322 631 324
rect 616 317 618 322
rect 629 317 631 322
rect 652 326 658 328
rect 652 324 654 326
rect 656 324 658 326
rect 652 322 658 324
rect 433 301 435 306
rect 440 301 442 306
rect 453 304 455 308
rect 481 305 483 310
rect 507 304 509 308
rect 520 301 522 306
rect 527 301 529 306
rect 560 301 562 306
rect 567 301 569 306
rect 580 304 582 308
rect 652 312 654 322
rect 663 321 665 336
rect 663 319 669 321
rect 663 317 665 319
rect 667 317 669 319
rect 659 315 669 317
rect 659 312 661 315
rect 609 301 611 306
rect 616 301 618 306
rect 629 304 631 308
rect 652 295 654 300
rect 659 295 661 300
rect 41 289 66 291
rect 41 281 43 289
rect 54 281 56 285
rect 64 281 66 289
rect 74 284 76 289
rect 81 284 83 289
rect 38 279 43 281
rect 38 276 40 279
rect 111 282 113 287
rect 121 282 123 287
rect 131 286 133 291
rect 54 269 56 272
rect 47 267 56 269
rect 64 268 66 272
rect 74 269 76 272
rect 38 259 40 267
rect 47 265 49 267
rect 51 265 56 267
rect 47 263 56 265
rect 72 267 76 269
rect 72 264 74 267
rect 54 259 56 263
rect 68 262 74 264
rect 81 263 83 272
rect 142 278 144 282
rect 166 280 168 285
rect 173 280 175 285
rect 213 289 238 291
rect 186 278 188 282
rect 213 281 215 289
rect 226 281 228 285
rect 236 281 238 289
rect 246 284 248 289
rect 253 284 255 289
rect 210 279 215 281
rect 210 276 212 279
rect 111 264 113 267
rect 121 264 123 267
rect 68 260 70 262
rect 72 260 74 262
rect 35 257 48 259
rect 54 257 64 259
rect 68 258 74 260
rect 35 256 37 257
rect 31 254 37 256
rect 46 254 48 257
rect 62 254 64 257
rect 72 254 74 258
rect 78 261 84 263
rect 78 259 80 261
rect 82 259 84 261
rect 78 257 84 259
rect 106 262 123 264
rect 106 260 108 262
rect 110 260 123 262
rect 106 258 123 260
rect 82 254 84 257
rect 111 254 113 258
rect 121 254 123 258
rect 131 264 133 267
rect 142 264 144 267
rect 131 262 144 264
rect 131 260 140 262
rect 142 260 144 262
rect 131 258 144 260
rect 131 254 133 258
rect 141 254 143 258
rect 166 256 168 269
rect 173 264 175 269
rect 186 264 188 269
rect 278 276 280 281
rect 457 278 459 282
rect 470 280 472 285
rect 477 280 479 285
rect 504 289 529 291
rect 504 281 506 289
rect 517 281 519 285
rect 527 281 529 289
rect 537 284 539 289
rect 544 284 546 289
rect 226 269 228 272
rect 219 267 228 269
rect 236 268 238 272
rect 246 269 248 272
rect 172 262 178 264
rect 172 260 174 262
rect 176 260 178 262
rect 172 258 178 260
rect 182 262 188 264
rect 182 260 184 262
rect 186 260 188 262
rect 182 258 188 260
rect 210 259 212 267
rect 219 265 221 267
rect 223 265 228 267
rect 219 263 228 265
rect 244 267 248 269
rect 244 264 246 267
rect 226 259 228 263
rect 240 262 246 264
rect 253 263 255 272
rect 501 279 506 281
rect 501 276 503 279
rect 278 264 280 267
rect 457 264 459 269
rect 470 264 472 269
rect 240 260 242 262
rect 244 260 246 262
rect 162 254 168 256
rect 31 252 33 254
rect 35 252 37 254
rect 31 250 37 252
rect 62 232 64 236
rect 72 232 74 236
rect 46 223 48 227
rect 162 252 164 254
rect 166 252 168 254
rect 162 250 168 252
rect 166 247 168 250
rect 176 247 178 258
rect 186 254 188 258
rect 207 257 220 259
rect 226 257 236 259
rect 240 258 246 260
rect 207 256 209 257
rect 203 254 209 256
rect 218 254 220 257
rect 234 254 236 257
rect 244 254 246 258
rect 250 261 256 263
rect 250 259 252 261
rect 254 259 256 261
rect 250 257 256 259
rect 254 254 256 257
rect 278 262 284 264
rect 278 260 280 262
rect 282 260 284 262
rect 278 258 284 260
rect 457 262 463 264
rect 457 260 459 262
rect 461 260 463 262
rect 457 258 463 260
rect 467 262 473 264
rect 467 260 469 262
rect 471 260 473 262
rect 467 258 473 260
rect 278 255 280 258
rect 111 231 113 236
rect 121 231 123 236
rect 131 231 133 236
rect 141 232 143 236
rect 203 252 205 254
rect 207 252 209 254
rect 203 250 209 252
rect 166 229 168 234
rect 176 229 178 234
rect 186 232 188 236
rect 82 223 84 227
rect 234 232 236 236
rect 244 232 246 236
rect 218 223 220 227
rect 457 254 459 258
rect 278 232 280 237
rect 467 247 469 258
rect 477 256 479 269
rect 581 280 583 285
rect 588 280 590 285
rect 517 269 519 272
rect 510 267 519 269
rect 527 268 529 272
rect 537 269 539 272
rect 501 259 503 267
rect 510 265 512 267
rect 514 265 519 267
rect 510 263 519 265
rect 535 267 539 269
rect 535 264 537 267
rect 517 259 519 263
rect 531 262 537 264
rect 544 263 546 272
rect 601 278 603 282
rect 629 276 631 281
rect 653 278 655 282
rect 664 281 666 286
rect 531 260 533 262
rect 535 260 537 262
rect 498 257 511 259
rect 517 257 527 259
rect 531 258 537 260
rect 498 256 500 257
rect 477 254 483 256
rect 477 252 479 254
rect 481 252 483 254
rect 477 250 483 252
rect 494 254 500 256
rect 509 254 511 257
rect 525 254 527 257
rect 535 254 537 258
rect 541 261 547 263
rect 541 259 543 261
rect 545 259 547 261
rect 541 257 547 259
rect 545 254 547 257
rect 581 256 583 269
rect 588 264 590 269
rect 601 264 603 269
rect 653 267 655 270
rect 629 264 631 267
rect 587 262 593 264
rect 587 260 589 262
rect 591 260 593 262
rect 587 258 593 260
rect 597 262 603 264
rect 597 260 599 262
rect 601 260 603 262
rect 597 258 603 260
rect 625 262 631 264
rect 625 260 627 262
rect 629 260 631 262
rect 651 265 657 267
rect 651 263 653 265
rect 655 263 657 265
rect 664 264 666 273
rect 651 261 657 263
rect 625 258 631 260
rect 577 254 583 256
rect 494 252 496 254
rect 498 252 500 254
rect 494 250 500 252
rect 477 247 479 250
rect 457 232 459 236
rect 254 223 256 227
rect 467 229 469 234
rect 477 229 479 234
rect 525 232 527 236
rect 535 232 537 236
rect 509 223 511 227
rect 577 252 579 254
rect 581 252 583 254
rect 577 250 583 252
rect 581 247 583 250
rect 591 247 593 258
rect 601 254 603 258
rect 629 255 631 258
rect 655 255 657 261
rect 661 262 667 264
rect 661 260 663 262
rect 665 260 667 262
rect 661 258 667 260
rect 662 255 664 258
rect 581 229 583 234
rect 591 229 593 234
rect 601 232 603 236
rect 629 232 631 237
rect 545 223 547 227
rect 655 223 657 227
rect 662 223 664 227
rect 38 215 40 219
rect 45 215 47 219
rect 55 215 57 219
rect 62 215 64 219
rect 162 215 164 219
rect 169 215 171 219
rect 179 215 181 219
rect 186 215 188 219
rect 92 205 94 210
rect 118 206 120 210
rect 128 208 130 213
rect 138 208 140 213
rect 38 179 40 188
rect 45 185 47 188
rect 55 185 57 188
rect 45 183 57 185
rect 50 182 57 183
rect 50 180 53 182
rect 55 180 57 182
rect 38 177 46 179
rect 38 176 42 177
rect 40 175 42 176
rect 44 175 46 177
rect 40 173 46 175
rect 50 178 57 180
rect 40 170 42 173
rect 50 170 52 178
rect 62 176 64 188
rect 92 184 94 187
rect 88 182 94 184
rect 88 180 90 182
rect 92 180 94 182
rect 88 178 94 180
rect 62 174 68 176
rect 92 175 94 178
rect 118 184 120 188
rect 128 184 130 195
rect 138 192 140 195
rect 138 190 144 192
rect 138 188 140 190
rect 142 188 144 190
rect 453 207 455 212
rect 463 207 465 212
rect 473 207 475 212
rect 515 215 517 219
rect 522 215 524 219
rect 529 215 531 219
rect 539 215 541 219
rect 546 215 548 219
rect 553 215 555 219
rect 587 215 589 219
rect 597 215 599 219
rect 621 215 623 219
rect 485 206 487 211
rect 138 186 144 188
rect 118 182 124 184
rect 118 180 120 182
rect 122 180 124 182
rect 118 178 124 180
rect 128 182 134 184
rect 128 180 130 182
rect 132 180 134 182
rect 128 178 134 180
rect 62 172 64 174
rect 66 172 68 174
rect 62 170 68 172
rect 118 173 120 178
rect 131 173 133 178
rect 138 173 140 186
rect 162 179 164 188
rect 169 185 171 188
rect 179 185 181 188
rect 169 183 181 185
rect 174 182 181 183
rect 174 180 177 182
rect 179 180 181 182
rect 162 177 170 179
rect 162 176 166 177
rect 164 175 166 176
rect 168 175 170 177
rect 164 173 170 175
rect 174 178 181 180
rect 92 161 94 166
rect 118 160 120 164
rect 164 170 166 173
rect 174 170 176 178
rect 186 176 188 188
rect 453 184 455 189
rect 463 184 465 194
rect 473 191 475 194
rect 473 189 479 191
rect 473 187 475 189
rect 477 187 479 189
rect 473 185 479 187
rect 453 182 459 184
rect 453 180 455 182
rect 457 180 459 182
rect 453 178 459 180
rect 463 182 469 184
rect 463 180 465 182
rect 467 180 469 182
rect 463 178 469 180
rect 186 174 192 176
rect 453 174 455 178
rect 466 174 468 178
rect 473 174 475 185
rect 485 184 487 193
rect 587 188 589 191
rect 485 182 491 184
rect 485 180 487 182
rect 489 180 491 182
rect 480 178 491 180
rect 480 174 482 178
rect 515 176 517 187
rect 522 184 524 187
rect 529 184 531 187
rect 539 184 541 187
rect 522 181 525 184
rect 529 182 541 184
rect 523 176 525 181
rect 539 176 541 182
rect 513 174 519 176
rect 186 172 188 174
rect 190 172 192 174
rect 186 170 192 172
rect 40 151 42 155
rect 50 151 52 155
rect 131 157 133 162
rect 138 157 140 162
rect 453 160 455 165
rect 513 172 515 174
rect 517 172 519 174
rect 513 170 519 172
rect 523 174 529 176
rect 523 172 525 174
rect 527 172 529 174
rect 523 170 529 172
rect 535 174 541 176
rect 535 172 537 174
rect 539 172 541 174
rect 546 178 548 187
rect 553 184 555 187
rect 578 186 589 188
rect 578 184 580 186
rect 582 184 589 186
rect 597 184 599 191
rect 657 215 659 219
rect 631 206 633 210
rect 641 206 643 210
rect 668 190 674 192
rect 668 188 670 190
rect 672 188 674 190
rect 553 182 562 184
rect 578 182 589 184
rect 556 180 558 182
rect 560 180 562 182
rect 556 178 562 180
rect 546 176 552 178
rect 546 174 548 176
rect 550 174 552 176
rect 587 175 589 182
rect 593 182 599 184
rect 593 180 595 182
rect 597 180 599 182
rect 593 178 599 180
rect 621 185 623 188
rect 621 183 627 185
rect 621 181 623 183
rect 625 181 627 183
rect 621 179 627 181
rect 631 184 633 188
rect 641 185 643 188
rect 657 185 659 188
rect 668 186 674 188
rect 668 185 670 186
rect 631 182 637 184
rect 641 183 651 185
rect 657 183 670 185
rect 631 180 633 182
rect 635 180 637 182
rect 594 175 596 178
rect 546 172 552 174
rect 535 170 541 172
rect 513 167 515 170
rect 525 167 527 170
rect 535 167 537 170
rect 164 151 166 155
rect 174 151 176 155
rect 466 156 468 161
rect 473 156 475 161
rect 480 156 482 161
rect 513 152 515 157
rect 525 152 527 157
rect 535 152 537 157
rect 622 170 624 179
rect 631 178 637 180
rect 649 179 651 183
rect 631 175 633 178
rect 629 173 633 175
rect 649 177 658 179
rect 649 175 654 177
rect 656 175 658 177
rect 665 175 667 183
rect 629 170 631 173
rect 639 170 641 174
rect 649 173 658 175
rect 649 170 651 173
rect 665 163 667 166
rect 662 161 667 163
rect 587 151 589 155
rect 594 151 596 155
rect 622 153 624 158
rect 629 153 631 158
rect 639 153 641 161
rect 649 157 651 161
rect 662 153 664 161
rect 639 151 664 153
rect 41 145 66 147
rect 41 137 43 145
rect 54 137 56 141
rect 64 137 66 145
rect 74 140 76 145
rect 81 140 83 145
rect 109 143 111 147
rect 116 143 118 147
rect 38 135 43 137
rect 38 132 40 135
rect 54 125 56 128
rect 47 123 56 125
rect 64 124 66 128
rect 74 125 76 128
rect 38 115 40 123
rect 47 121 49 123
rect 51 121 56 123
rect 47 119 56 121
rect 72 123 76 125
rect 72 120 74 123
rect 54 115 56 119
rect 68 118 74 120
rect 81 119 83 128
rect 144 136 146 141
rect 151 136 153 141
rect 164 134 166 138
rect 192 132 194 137
rect 109 120 111 123
rect 68 116 70 118
rect 72 116 74 118
rect 35 113 48 115
rect 54 113 64 115
rect 68 114 74 116
rect 35 112 37 113
rect 31 110 37 112
rect 46 110 48 113
rect 62 110 64 113
rect 72 110 74 114
rect 78 117 84 119
rect 78 115 80 117
rect 82 115 84 117
rect 78 113 84 115
rect 82 110 84 113
rect 106 118 112 120
rect 106 116 108 118
rect 110 116 112 118
rect 106 114 112 116
rect 116 116 118 123
rect 116 114 127 116
rect 31 108 33 110
rect 35 108 37 110
rect 31 106 37 108
rect 62 88 64 92
rect 72 88 74 92
rect 46 79 48 83
rect 106 107 108 114
rect 116 112 123 114
rect 125 112 127 114
rect 144 112 146 125
rect 151 120 153 125
rect 164 120 166 125
rect 441 140 459 142
rect 441 136 443 140
rect 457 137 459 140
rect 467 137 469 142
rect 479 137 481 142
rect 489 137 491 142
rect 530 137 532 142
rect 537 137 539 142
rect 544 137 546 142
rect 437 134 443 136
rect 437 132 439 134
rect 441 132 443 134
rect 437 130 443 132
rect 447 126 453 128
rect 437 123 443 125
rect 150 118 156 120
rect 150 116 152 118
rect 154 116 156 118
rect 150 114 156 116
rect 160 118 166 120
rect 160 116 162 118
rect 164 116 166 118
rect 160 114 166 116
rect 116 110 127 112
rect 140 110 146 112
rect 116 107 118 110
rect 140 108 142 110
rect 144 108 146 110
rect 140 106 146 108
rect 144 103 146 106
rect 154 103 156 114
rect 164 110 166 114
rect 192 120 194 123
rect 437 121 439 123
rect 441 121 443 123
rect 192 118 198 120
rect 437 119 443 121
rect 447 124 449 126
rect 451 124 453 126
rect 447 122 453 124
rect 192 116 194 118
rect 196 116 198 118
rect 192 114 198 116
rect 427 117 433 119
rect 427 115 429 117
rect 431 115 433 117
rect 192 111 194 114
rect 427 113 435 115
rect 433 110 435 113
rect 440 110 442 119
rect 447 110 449 122
rect 457 115 459 131
rect 467 128 469 131
rect 466 126 472 128
rect 479 126 481 131
rect 466 124 468 126
rect 470 124 472 126
rect 466 122 472 124
rect 470 116 472 122
rect 477 124 483 126
rect 477 122 479 124
rect 481 122 483 124
rect 477 120 483 122
rect 454 113 466 115
rect 470 113 473 116
rect 454 110 456 113
rect 464 110 466 113
rect 471 110 473 113
rect 478 110 480 120
rect 489 119 491 131
rect 557 133 559 138
rect 581 136 583 141
rect 588 136 590 141
rect 655 143 657 147
rect 662 143 664 147
rect 601 134 603 138
rect 629 132 631 137
rect 530 120 532 124
rect 489 117 498 119
rect 489 115 494 117
rect 496 115 498 117
rect 485 113 498 115
rect 521 118 532 120
rect 521 116 523 118
rect 525 116 527 118
rect 521 114 527 116
rect 485 110 487 113
rect 144 85 146 90
rect 154 85 156 90
rect 164 88 166 92
rect 192 88 194 93
rect 433 88 435 92
rect 440 88 442 92
rect 447 88 449 92
rect 454 88 456 92
rect 82 79 84 83
rect 106 79 108 83
rect 116 79 118 83
rect 525 105 527 114
rect 537 113 539 124
rect 544 120 546 124
rect 557 120 559 124
rect 543 118 549 120
rect 543 116 545 118
rect 547 116 549 118
rect 543 114 549 116
rect 553 118 559 120
rect 553 116 555 118
rect 557 116 559 118
rect 553 114 559 116
rect 533 111 539 113
rect 533 109 535 111
rect 537 109 539 111
rect 533 107 539 109
rect 537 104 539 107
rect 547 104 549 114
rect 557 109 559 114
rect 581 112 583 125
rect 588 120 590 125
rect 601 120 603 125
rect 629 120 631 123
rect 587 118 593 120
rect 587 116 589 118
rect 591 116 593 118
rect 587 114 593 116
rect 597 118 603 120
rect 597 116 599 118
rect 601 116 603 118
rect 597 114 603 116
rect 625 118 631 120
rect 625 116 627 118
rect 629 116 631 118
rect 655 116 657 123
rect 662 120 664 123
rect 625 114 631 116
rect 577 110 583 112
rect 525 87 527 92
rect 577 108 579 110
rect 581 108 583 110
rect 577 106 583 108
rect 581 103 583 106
rect 591 103 593 114
rect 601 110 603 114
rect 629 111 631 114
rect 646 114 657 116
rect 661 118 667 120
rect 661 116 663 118
rect 665 116 667 118
rect 661 114 667 116
rect 646 112 648 114
rect 650 112 657 114
rect 464 80 466 85
rect 471 80 473 85
rect 478 80 480 85
rect 485 80 487 85
rect 537 86 539 91
rect 547 86 549 91
rect 557 86 559 91
rect 646 110 657 112
rect 655 107 657 110
rect 665 107 667 114
rect 581 85 583 90
rect 591 85 593 90
rect 601 88 603 92
rect 629 88 631 93
rect 655 79 657 83
rect 665 79 667 83
rect 38 71 40 75
rect 45 71 47 75
rect 55 71 57 75
rect 62 71 64 75
rect 117 71 119 75
rect 90 61 92 66
rect 38 35 40 44
rect 45 41 47 44
rect 55 41 57 44
rect 45 39 57 41
rect 50 38 57 39
rect 50 36 53 38
rect 55 36 57 38
rect 38 33 46 35
rect 38 32 42 33
rect 40 31 42 32
rect 44 31 46 33
rect 40 29 46 31
rect 50 34 57 36
rect 40 26 42 29
rect 50 26 52 34
rect 62 32 64 44
rect 153 71 155 75
rect 127 62 129 66
rect 137 62 139 66
rect 198 70 200 74
rect 188 62 190 66
rect 164 46 170 48
rect 417 67 419 72
rect 427 67 429 72
rect 437 67 439 72
rect 447 67 449 72
rect 473 71 475 75
rect 387 61 389 66
rect 164 44 166 46
rect 168 44 170 46
rect 90 40 92 43
rect 86 38 92 40
rect 86 36 88 38
rect 90 36 92 38
rect 86 34 92 36
rect 117 41 119 44
rect 117 39 123 41
rect 117 37 119 39
rect 121 37 123 39
rect 117 35 123 37
rect 127 40 129 44
rect 137 41 139 44
rect 153 41 155 44
rect 164 42 170 44
rect 164 41 166 42
rect 188 41 190 46
rect 198 41 200 46
rect 127 38 133 40
rect 137 39 147 41
rect 153 39 166 41
rect 180 39 200 41
rect 387 40 389 43
rect 417 40 419 50
rect 427 47 429 50
rect 437 47 439 50
rect 423 45 429 47
rect 423 43 425 45
rect 427 43 429 45
rect 423 41 429 43
rect 433 45 439 47
rect 433 43 435 45
rect 437 43 439 45
rect 433 41 439 43
rect 127 36 129 38
rect 131 36 133 38
rect 62 30 68 32
rect 90 31 92 34
rect 62 28 64 30
rect 66 28 68 30
rect 62 26 68 28
rect 118 26 120 35
rect 127 34 133 36
rect 145 35 147 39
rect 127 31 129 34
rect 125 29 129 31
rect 145 33 154 35
rect 145 31 150 33
rect 152 31 154 33
rect 161 31 163 39
rect 180 37 182 39
rect 184 37 190 39
rect 180 35 190 37
rect 188 31 190 35
rect 198 31 200 39
rect 383 38 389 40
rect 383 36 385 38
rect 387 36 389 38
rect 383 34 389 36
rect 411 38 419 40
rect 411 36 413 38
rect 415 36 419 38
rect 411 34 422 36
rect 387 31 389 34
rect 420 31 422 34
rect 427 31 429 41
rect 434 31 436 41
rect 447 40 449 50
rect 509 71 511 75
rect 483 62 485 66
rect 493 62 495 66
rect 587 71 589 75
rect 594 71 596 75
rect 621 71 623 75
rect 541 64 543 69
rect 551 64 553 69
rect 561 62 563 66
rect 541 48 543 51
rect 520 46 526 48
rect 520 44 522 46
rect 524 44 526 46
rect 443 38 449 40
rect 443 37 445 38
rect 441 36 445 37
rect 447 36 449 38
rect 441 34 449 36
rect 473 41 475 44
rect 473 39 479 41
rect 473 37 475 39
rect 477 37 479 39
rect 473 35 479 37
rect 483 40 485 44
rect 493 41 495 44
rect 509 41 511 44
rect 520 42 526 44
rect 537 46 543 48
rect 537 44 539 46
rect 541 44 543 46
rect 537 42 543 44
rect 520 41 522 42
rect 483 38 489 40
rect 493 39 503 41
rect 509 39 522 41
rect 483 36 485 38
rect 487 36 489 38
rect 441 31 443 34
rect 125 26 127 29
rect 135 26 137 30
rect 145 29 154 31
rect 145 26 147 29
rect 90 17 92 22
rect 161 19 163 22
rect 158 17 163 19
rect 40 7 42 11
rect 50 7 52 11
rect 118 9 120 14
rect 125 9 127 14
rect 135 9 137 17
rect 145 13 147 17
rect 158 9 160 17
rect 188 16 190 21
rect 198 16 200 21
rect 387 17 389 22
rect 135 7 160 9
rect 474 26 476 35
rect 483 34 489 36
rect 501 35 503 39
rect 483 31 485 34
rect 481 29 485 31
rect 501 33 510 35
rect 501 31 506 33
rect 508 31 510 33
rect 517 31 519 39
rect 481 26 483 29
rect 491 26 493 30
rect 501 29 510 31
rect 501 26 503 29
rect 541 29 543 42
rect 551 40 553 51
rect 561 40 563 44
rect 657 71 659 75
rect 631 62 633 66
rect 641 62 643 66
rect 668 46 674 48
rect 668 44 670 46
rect 672 44 674 46
rect 547 38 553 40
rect 547 36 549 38
rect 551 36 553 38
rect 547 34 553 36
rect 557 38 563 40
rect 557 36 559 38
rect 561 36 563 38
rect 587 37 589 43
rect 594 40 596 43
rect 621 41 623 44
rect 557 34 563 36
rect 548 29 550 34
rect 561 29 563 34
rect 583 35 589 37
rect 583 33 585 35
rect 587 33 589 35
rect 593 38 599 40
rect 593 36 595 38
rect 597 36 599 38
rect 593 34 599 36
rect 621 39 627 41
rect 621 37 623 39
rect 625 37 627 39
rect 621 35 627 37
rect 631 40 633 44
rect 641 41 643 44
rect 657 41 659 44
rect 668 42 674 44
rect 668 41 670 42
rect 631 38 637 40
rect 641 39 651 41
rect 657 39 670 41
rect 631 36 633 38
rect 635 36 637 38
rect 583 31 589 33
rect 517 19 519 22
rect 514 17 519 19
rect 585 28 587 31
rect 596 25 598 34
rect 622 26 624 35
rect 631 34 637 36
rect 649 35 651 39
rect 631 31 633 34
rect 629 29 633 31
rect 649 33 658 35
rect 649 31 654 33
rect 656 31 658 33
rect 665 31 667 39
rect 629 26 631 29
rect 639 26 641 30
rect 649 29 658 31
rect 649 26 651 29
rect 420 7 422 11
rect 427 7 429 11
rect 434 7 436 11
rect 441 7 443 11
rect 474 9 476 14
rect 481 9 483 14
rect 491 9 493 17
rect 501 13 503 17
rect 514 9 516 17
rect 491 7 516 9
rect 541 13 543 18
rect 548 13 550 18
rect 561 16 563 20
rect 585 16 587 20
rect 596 12 598 17
rect 665 19 667 22
rect 662 17 667 19
rect 622 9 624 14
rect 629 9 631 14
rect 639 9 641 17
rect 649 13 651 17
rect 662 9 664 17
rect 639 7 664 9
<< ndif >>
rect 85 720 91 722
rect 85 718 87 720
rect 89 718 91 720
rect 85 716 91 718
rect 69 713 74 716
rect 45 711 54 713
rect 45 709 47 711
rect 49 709 54 711
rect 45 708 54 709
rect 33 705 38 708
rect 31 703 38 705
rect 31 701 33 703
rect 35 701 38 703
rect 31 699 38 701
rect 40 704 54 708
rect 56 708 64 713
rect 56 706 59 708
rect 61 706 64 708
rect 56 704 64 706
rect 66 710 74 713
rect 66 708 69 710
rect 71 708 74 710
rect 66 704 74 708
rect 76 704 81 716
rect 83 704 91 716
rect 99 720 105 722
rect 99 718 101 720
rect 103 718 105 720
rect 99 713 105 718
rect 146 720 153 722
rect 146 718 148 720
rect 150 718 153 720
rect 99 705 107 713
rect 109 711 116 713
rect 109 709 112 711
rect 114 710 116 711
rect 146 712 153 718
rect 233 720 239 722
rect 233 718 235 720
rect 237 718 239 720
rect 287 720 294 722
rect 287 719 289 720
rect 233 716 239 718
rect 217 713 222 716
rect 146 710 155 712
rect 114 709 118 710
rect 109 705 118 709
rect 40 699 45 704
rect 113 702 118 705
rect 120 708 127 710
rect 120 706 123 708
rect 125 706 127 708
rect 120 702 127 706
rect 135 708 142 710
rect 135 706 137 708
rect 139 706 142 708
rect 135 704 142 706
rect 137 701 142 704
rect 144 701 155 710
rect 157 701 162 712
rect 164 710 171 712
rect 164 708 167 710
rect 169 708 171 710
rect 193 711 202 713
rect 193 709 195 711
rect 197 709 202 711
rect 193 708 202 709
rect 164 706 171 708
rect 164 701 169 706
rect 181 705 186 708
rect 179 703 186 705
rect 179 701 181 703
rect 183 701 186 703
rect 179 699 186 701
rect 188 704 202 708
rect 204 708 212 713
rect 204 706 207 708
rect 209 706 212 708
rect 204 704 212 706
rect 214 710 222 713
rect 214 708 217 710
rect 219 708 222 710
rect 214 704 222 708
rect 224 704 229 716
rect 231 704 239 716
rect 257 713 262 719
rect 255 711 262 713
rect 255 709 257 711
rect 259 709 262 711
rect 255 707 262 709
rect 188 699 193 704
rect 257 699 262 707
rect 264 699 269 719
rect 271 699 276 719
rect 278 699 283 719
rect 285 718 289 719
rect 291 718 294 720
rect 285 699 294 718
rect 497 710 503 712
rect 497 708 499 710
rect 501 709 503 710
rect 589 720 595 722
rect 589 718 591 720
rect 593 718 595 720
rect 589 716 595 718
rect 573 713 578 716
rect 549 711 558 713
rect 501 708 505 709
rect 311 705 316 708
rect 309 703 316 705
rect 309 701 311 703
rect 313 701 316 703
rect 309 699 316 701
rect 318 706 329 708
rect 318 704 325 706
rect 327 704 329 706
rect 318 699 329 704
rect 497 699 505 708
rect 507 703 515 709
rect 507 701 510 703
rect 512 701 515 703
rect 507 699 515 701
rect 517 707 525 709
rect 549 709 551 711
rect 553 709 558 711
rect 549 708 558 709
rect 517 705 521 707
rect 523 705 525 707
rect 537 705 542 708
rect 517 699 525 705
rect 535 703 542 705
rect 535 701 537 703
rect 539 701 542 703
rect 535 699 542 701
rect 544 704 558 708
rect 560 708 568 713
rect 560 706 563 708
rect 565 706 568 708
rect 560 704 568 706
rect 570 710 578 713
rect 570 708 573 710
rect 575 708 578 710
rect 570 704 578 708
rect 580 704 585 716
rect 587 704 595 716
rect 608 705 613 708
rect 544 699 549 704
rect 606 703 613 705
rect 606 701 608 703
rect 610 701 613 703
rect 606 699 613 701
rect 615 706 626 708
rect 645 717 653 719
rect 645 715 648 717
rect 650 715 653 717
rect 645 710 653 715
rect 645 708 648 710
rect 650 708 653 710
rect 615 704 622 706
rect 624 704 626 706
rect 645 704 653 708
rect 655 710 663 719
rect 655 708 658 710
rect 660 708 663 710
rect 655 704 663 708
rect 665 717 673 719
rect 665 715 668 717
rect 670 715 673 717
rect 665 704 673 715
rect 615 699 626 704
rect 36 599 41 607
rect 34 597 41 599
rect 34 595 36 597
rect 38 595 41 597
rect 34 593 41 595
rect 36 587 41 593
rect 43 587 48 607
rect 50 598 59 607
rect 67 605 74 607
rect 67 603 69 605
rect 71 603 74 605
rect 67 601 74 603
rect 69 598 74 601
rect 76 602 87 607
rect 97 602 102 605
rect 76 600 83 602
rect 85 600 87 602
rect 76 598 87 600
rect 95 600 102 602
rect 95 598 97 600
rect 99 598 102 600
rect 50 596 55 598
rect 57 596 59 598
rect 50 591 59 596
rect 95 596 102 598
rect 104 596 115 605
rect 106 594 115 596
rect 117 594 122 605
rect 124 600 129 605
rect 139 604 146 606
rect 139 602 141 604
rect 143 602 146 604
rect 139 600 146 602
rect 124 598 131 600
rect 124 596 127 598
rect 129 596 131 598
rect 141 597 146 600
rect 148 597 159 606
rect 124 594 131 596
rect 50 589 55 591
rect 57 589 59 591
rect 50 587 59 589
rect 106 588 113 594
rect 150 593 159 597
rect 161 593 166 606
rect 168 593 173 606
rect 175 599 180 606
rect 175 597 182 599
rect 175 595 178 597
rect 180 595 182 597
rect 175 593 182 595
rect 207 597 214 599
rect 207 595 209 597
rect 211 595 214 597
rect 207 593 214 595
rect 216 597 224 599
rect 216 595 219 597
rect 221 595 224 597
rect 216 593 224 595
rect 226 593 236 599
rect 238 597 246 599
rect 238 595 241 597
rect 243 595 246 597
rect 238 593 246 595
rect 248 597 255 599
rect 248 595 251 597
rect 253 595 255 597
rect 248 593 255 595
rect 106 586 108 588
rect 110 586 113 588
rect 106 584 113 586
rect 150 588 157 593
rect 228 588 234 593
rect 500 602 511 607
rect 500 600 502 602
rect 504 600 511 602
rect 500 598 511 600
rect 513 605 520 607
rect 513 603 516 605
rect 518 603 520 605
rect 513 601 520 603
rect 534 602 539 605
rect 513 598 518 601
rect 532 600 539 602
rect 532 598 534 600
rect 536 598 539 600
rect 532 596 539 598
rect 541 596 552 605
rect 543 594 552 596
rect 554 594 559 605
rect 561 600 566 605
rect 561 598 568 600
rect 561 596 564 598
rect 566 596 568 598
rect 561 594 568 596
rect 578 598 587 607
rect 578 596 580 598
rect 582 596 587 598
rect 150 586 152 588
rect 154 586 157 588
rect 150 584 157 586
rect 228 586 230 588
rect 232 586 234 588
rect 228 584 234 586
rect 543 588 550 594
rect 578 591 587 596
rect 578 589 580 591
rect 582 589 587 591
rect 543 586 545 588
rect 547 586 550 588
rect 578 587 587 589
rect 589 587 594 607
rect 596 599 601 607
rect 660 602 665 607
rect 596 597 603 599
rect 596 595 599 597
rect 601 595 603 597
rect 596 593 603 595
rect 596 587 601 593
rect 614 590 622 602
rect 624 590 629 602
rect 631 598 639 602
rect 631 596 634 598
rect 636 596 639 598
rect 631 593 639 596
rect 641 600 649 602
rect 641 598 644 600
rect 646 598 649 600
rect 641 593 649 598
rect 651 598 665 602
rect 667 605 674 607
rect 667 603 670 605
rect 672 603 674 605
rect 667 601 674 603
rect 667 598 672 601
rect 651 597 660 598
rect 651 595 656 597
rect 658 595 660 597
rect 651 593 660 595
rect 631 590 636 593
rect 614 588 620 590
rect 543 584 550 586
rect 614 586 616 588
rect 618 586 620 588
rect 614 584 620 586
rect 85 576 91 578
rect 85 574 87 576
rect 89 574 91 576
rect 85 572 91 574
rect 69 569 74 572
rect 45 567 54 569
rect 45 565 47 567
rect 49 565 54 567
rect 45 564 54 565
rect 33 561 38 564
rect 31 559 38 561
rect 31 557 33 559
rect 35 557 38 559
rect 31 555 38 557
rect 40 560 54 564
rect 56 564 64 569
rect 56 562 59 564
rect 61 562 64 564
rect 56 560 64 562
rect 66 566 74 569
rect 66 564 69 566
rect 71 564 74 566
rect 66 560 74 564
rect 76 560 81 572
rect 83 560 91 572
rect 104 569 109 575
rect 102 567 109 569
rect 102 565 104 567
rect 106 565 109 567
rect 102 563 109 565
rect 40 555 45 560
rect 104 555 109 563
rect 111 555 116 575
rect 118 573 127 575
rect 118 571 123 573
rect 125 571 127 573
rect 118 566 127 571
rect 118 564 123 566
rect 125 564 127 566
rect 118 555 127 564
rect 159 576 166 578
rect 159 574 162 576
rect 164 574 166 576
rect 159 573 166 574
rect 182 576 188 578
rect 182 574 184 576
rect 186 574 188 576
rect 182 573 188 574
rect 241 576 248 578
rect 241 574 244 576
rect 246 574 248 576
rect 159 563 168 573
rect 170 567 178 573
rect 170 565 173 567
rect 175 565 178 567
rect 170 563 178 565
rect 180 563 190 573
rect 192 569 197 573
rect 241 569 248 574
rect 576 576 583 578
rect 192 567 199 569
rect 192 565 195 567
rect 197 565 199 567
rect 192 563 199 565
rect 216 567 223 569
rect 216 565 218 567
rect 220 565 223 567
rect 216 563 223 565
rect 218 556 223 563
rect 225 556 230 569
rect 232 556 237 569
rect 239 565 248 569
rect 239 556 250 565
rect 252 562 257 565
rect 252 560 259 562
rect 444 561 449 564
rect 252 558 255 560
rect 257 558 259 560
rect 252 556 259 558
rect 442 559 449 561
rect 442 557 444 559
rect 446 557 449 559
rect 442 555 449 557
rect 451 562 462 564
rect 521 573 529 575
rect 521 571 524 573
rect 526 571 529 573
rect 521 566 529 571
rect 521 564 524 566
rect 526 564 529 566
rect 451 560 458 562
rect 460 560 462 562
rect 521 560 529 564
rect 531 566 539 575
rect 531 564 534 566
rect 536 564 539 566
rect 531 560 539 564
rect 541 573 549 575
rect 576 574 579 576
rect 581 574 583 576
rect 541 571 544 573
rect 546 571 549 573
rect 541 560 549 571
rect 576 568 583 574
rect 558 566 565 568
rect 558 564 560 566
rect 562 564 565 566
rect 558 562 565 564
rect 451 555 462 560
rect 560 557 565 562
rect 567 557 572 568
rect 574 566 583 568
rect 574 557 585 566
rect 587 564 594 566
rect 587 562 590 564
rect 592 562 594 564
rect 587 560 594 562
rect 606 561 611 564
rect 587 557 592 560
rect 604 559 611 561
rect 604 557 606 559
rect 608 557 611 559
rect 604 555 611 557
rect 613 562 624 564
rect 645 573 653 575
rect 645 571 648 573
rect 650 571 653 573
rect 645 566 653 571
rect 645 564 648 566
rect 650 564 653 566
rect 613 560 620 562
rect 622 560 624 562
rect 645 560 653 564
rect 655 566 663 575
rect 655 564 658 566
rect 660 564 663 566
rect 655 560 663 564
rect 665 573 673 575
rect 665 571 668 573
rect 670 571 673 573
rect 665 560 673 571
rect 613 555 624 560
rect 67 461 74 463
rect 45 457 50 460
rect 31 454 39 457
rect 28 450 39 454
rect 31 449 39 450
rect 41 453 50 457
rect 41 451 44 453
rect 46 452 50 453
rect 52 456 59 460
rect 67 459 69 461
rect 71 459 74 461
rect 67 457 74 459
rect 52 454 55 456
rect 57 454 59 456
rect 69 454 74 457
rect 76 458 87 463
rect 97 458 102 461
rect 76 456 83 458
rect 85 456 87 458
rect 76 454 87 456
rect 95 456 102 458
rect 95 454 97 456
rect 99 454 102 456
rect 52 452 59 454
rect 46 451 48 452
rect 41 449 48 451
rect 31 444 37 449
rect 95 452 102 454
rect 104 452 115 461
rect 106 450 115 452
rect 117 450 122 461
rect 124 456 129 461
rect 197 458 202 463
rect 124 454 131 456
rect 124 452 127 454
rect 129 452 131 454
rect 124 450 131 452
rect 31 442 33 444
rect 35 442 37 444
rect 31 440 37 442
rect 106 444 113 450
rect 151 446 159 458
rect 161 446 166 458
rect 168 454 176 458
rect 168 452 171 454
rect 173 452 176 454
rect 168 449 176 452
rect 178 456 186 458
rect 178 454 181 456
rect 183 454 186 456
rect 178 449 186 454
rect 188 454 202 458
rect 204 461 211 463
rect 204 459 207 461
rect 209 459 211 461
rect 204 457 211 459
rect 204 454 209 457
rect 221 456 226 461
rect 219 454 226 456
rect 188 453 197 454
rect 188 451 193 453
rect 195 451 197 453
rect 188 449 197 451
rect 219 452 221 454
rect 223 452 226 454
rect 219 450 226 452
rect 228 450 233 461
rect 235 452 246 461
rect 248 458 253 461
rect 488 458 493 463
rect 248 456 255 458
rect 248 454 251 456
rect 253 454 255 456
rect 248 452 255 454
rect 235 450 244 452
rect 168 446 173 449
rect 106 442 108 444
rect 110 442 113 444
rect 106 440 113 442
rect 151 444 157 446
rect 151 442 153 444
rect 155 442 157 444
rect 151 440 157 442
rect 237 444 244 450
rect 442 446 450 458
rect 452 446 457 458
rect 459 454 467 458
rect 459 452 462 454
rect 464 452 467 454
rect 459 449 467 452
rect 469 456 477 458
rect 469 454 472 456
rect 474 454 477 456
rect 469 449 477 454
rect 479 454 493 458
rect 495 461 502 463
rect 554 461 561 463
rect 495 459 498 461
rect 500 459 502 461
rect 495 457 502 459
rect 512 458 517 461
rect 495 454 500 457
rect 510 456 517 458
rect 510 454 512 456
rect 514 454 517 456
rect 479 453 488 454
rect 479 451 484 453
rect 486 451 488 453
rect 510 452 517 454
rect 519 452 530 461
rect 479 449 488 451
rect 459 446 464 449
rect 237 442 240 444
rect 242 442 244 444
rect 237 440 244 442
rect 442 444 448 446
rect 442 442 444 444
rect 446 442 448 444
rect 442 440 448 442
rect 521 450 530 452
rect 532 450 537 461
rect 539 456 544 461
rect 554 459 556 461
rect 558 459 561 461
rect 554 457 561 459
rect 539 454 546 456
rect 539 452 542 454
rect 544 452 546 454
rect 556 452 561 457
rect 563 452 572 463
rect 539 450 546 452
rect 521 444 528 450
rect 565 450 567 452
rect 569 450 572 452
rect 521 442 523 444
rect 525 442 528 444
rect 521 440 528 442
rect 565 444 572 450
rect 574 460 582 463
rect 574 458 577 460
rect 579 458 582 460
rect 574 453 582 458
rect 574 451 577 453
rect 579 451 582 453
rect 574 448 582 451
rect 584 461 592 463
rect 584 459 587 461
rect 589 459 592 461
rect 584 448 592 459
rect 594 455 599 463
rect 660 458 665 463
rect 594 453 601 455
rect 594 451 597 453
rect 599 451 601 453
rect 594 448 601 451
rect 574 444 579 448
rect 614 446 622 458
rect 624 446 629 458
rect 631 454 639 458
rect 631 452 634 454
rect 636 452 639 454
rect 631 449 639 452
rect 641 456 649 458
rect 641 454 644 456
rect 646 454 649 456
rect 641 449 649 454
rect 651 454 665 458
rect 667 461 674 463
rect 667 459 670 461
rect 672 459 674 461
rect 667 457 674 459
rect 667 454 672 457
rect 651 453 660 454
rect 651 451 656 453
rect 658 451 660 453
rect 651 449 660 451
rect 631 446 636 449
rect 614 444 620 446
rect 614 442 616 444
rect 618 442 620 444
rect 614 440 620 442
rect 32 428 44 430
rect 32 426 34 428
rect 36 426 44 428
rect 32 418 44 426
rect 46 418 51 430
rect 53 424 58 430
rect 78 432 85 434
rect 78 430 80 432
rect 82 430 85 432
rect 53 422 60 424
rect 78 424 85 430
rect 127 432 134 434
rect 127 430 129 432
rect 131 430 134 432
rect 78 422 87 424
rect 53 420 56 422
rect 58 420 60 422
rect 53 418 60 420
rect 67 420 74 422
rect 67 418 69 420
rect 71 418 74 420
rect 67 416 74 418
rect 69 413 74 416
rect 76 413 87 422
rect 89 413 94 424
rect 96 422 103 424
rect 127 424 134 430
rect 187 432 194 434
rect 187 430 190 432
rect 192 430 194 432
rect 187 424 194 430
rect 254 432 261 434
rect 254 430 256 432
rect 258 430 261 432
rect 127 422 136 424
rect 96 420 99 422
rect 101 420 103 422
rect 96 418 103 420
rect 116 420 123 422
rect 116 418 118 420
rect 120 418 123 420
rect 96 413 101 418
rect 116 416 123 418
rect 118 413 123 416
rect 125 413 136 422
rect 138 413 143 424
rect 145 422 152 424
rect 145 420 148 422
rect 150 420 152 422
rect 145 418 152 420
rect 169 422 176 424
rect 169 420 171 422
rect 173 420 176 422
rect 169 418 176 420
rect 145 413 150 418
rect 171 413 176 418
rect 178 413 183 424
rect 185 422 194 424
rect 185 413 196 422
rect 198 420 205 422
rect 254 424 261 430
rect 298 432 305 434
rect 298 430 300 432
rect 302 430 305 432
rect 435 432 442 434
rect 435 430 438 432
rect 440 430 442 432
rect 254 422 263 424
rect 243 420 250 422
rect 198 418 201 420
rect 203 418 205 420
rect 198 416 205 418
rect 217 417 222 420
rect 198 413 203 416
rect 215 415 222 417
rect 215 413 217 415
rect 219 413 222 415
rect 215 411 222 413
rect 224 418 235 420
rect 224 416 231 418
rect 233 416 235 418
rect 243 418 245 420
rect 247 418 250 420
rect 243 416 250 418
rect 224 411 235 416
rect 245 413 250 416
rect 252 413 263 422
rect 265 413 270 424
rect 272 422 279 424
rect 272 420 275 422
rect 277 420 279 422
rect 298 425 305 430
rect 298 421 307 425
rect 272 418 279 420
rect 289 418 294 421
rect 272 413 277 418
rect 287 416 294 418
rect 287 414 289 416
rect 291 414 294 416
rect 287 412 294 414
rect 296 412 307 421
rect 309 412 314 425
rect 316 412 321 425
rect 323 423 330 425
rect 435 424 442 430
rect 508 432 515 434
rect 508 430 511 432
rect 513 430 515 432
rect 323 421 326 423
rect 328 421 330 423
rect 323 419 330 421
rect 417 422 424 424
rect 417 420 419 422
rect 421 420 424 422
rect 323 412 328 419
rect 417 418 424 420
rect 419 413 424 418
rect 426 413 431 424
rect 433 422 442 424
rect 433 413 444 422
rect 446 420 453 422
rect 508 424 515 430
rect 549 432 556 434
rect 549 430 551 432
rect 553 430 556 432
rect 612 432 619 434
rect 612 430 615 432
rect 617 430 619 432
rect 490 422 497 424
rect 490 420 492 422
rect 494 420 497 422
rect 446 418 449 420
rect 451 418 453 420
rect 446 416 453 418
rect 464 417 469 420
rect 446 413 451 416
rect 462 415 469 417
rect 462 413 464 415
rect 466 413 469 415
rect 462 411 469 413
rect 471 418 482 420
rect 490 418 497 420
rect 471 416 478 418
rect 480 416 482 418
rect 471 411 482 416
rect 492 413 497 418
rect 499 413 504 424
rect 506 422 515 424
rect 549 424 556 430
rect 612 425 619 430
rect 640 431 646 433
rect 640 430 648 431
rect 640 428 642 430
rect 644 428 648 430
rect 549 422 558 424
rect 506 413 517 422
rect 519 420 526 422
rect 519 418 522 420
rect 524 418 526 420
rect 519 416 526 418
rect 538 420 545 422
rect 538 418 540 420
rect 542 418 545 420
rect 538 416 545 418
rect 519 413 524 416
rect 540 413 545 416
rect 547 413 558 422
rect 560 413 565 424
rect 567 422 574 424
rect 567 420 570 422
rect 572 420 574 422
rect 567 418 574 420
rect 587 423 594 425
rect 587 421 589 423
rect 591 421 594 423
rect 587 419 594 421
rect 567 413 572 418
rect 589 412 594 419
rect 596 412 601 425
rect 603 412 608 425
rect 610 421 619 425
rect 610 412 621 421
rect 623 418 628 421
rect 623 416 630 418
rect 623 414 626 416
rect 628 414 630 416
rect 623 412 630 414
rect 640 411 648 428
rect 650 411 655 431
rect 657 411 662 431
rect 664 425 669 431
rect 664 423 671 425
rect 664 421 667 423
rect 669 421 671 423
rect 664 419 671 421
rect 664 411 669 419
rect 36 311 41 319
rect 34 309 41 311
rect 34 307 36 309
rect 38 307 41 309
rect 34 305 41 307
rect 36 299 41 305
rect 43 299 48 319
rect 50 299 55 319
rect 57 302 65 319
rect 75 316 82 318
rect 75 314 77 316
rect 79 314 82 316
rect 75 312 82 314
rect 77 309 82 312
rect 84 309 95 318
rect 86 305 95 309
rect 97 305 102 318
rect 104 305 109 318
rect 111 311 116 318
rect 133 312 138 317
rect 111 309 118 311
rect 111 307 114 309
rect 116 307 118 309
rect 111 305 118 307
rect 131 310 138 312
rect 131 308 133 310
rect 135 308 138 310
rect 131 306 138 308
rect 140 306 145 317
rect 147 308 158 317
rect 160 314 165 317
rect 181 314 186 317
rect 160 312 167 314
rect 160 310 163 312
rect 165 310 167 312
rect 160 308 167 310
rect 179 312 186 314
rect 179 310 181 312
rect 183 310 186 312
rect 179 308 186 310
rect 188 308 199 317
rect 147 306 156 308
rect 57 300 61 302
rect 63 300 65 302
rect 57 299 65 300
rect 59 297 65 299
rect 86 300 93 305
rect 149 300 156 306
rect 190 306 199 308
rect 201 306 206 317
rect 208 312 213 317
rect 223 314 234 319
rect 223 312 225 314
rect 227 312 234 314
rect 208 310 215 312
rect 223 310 234 312
rect 236 317 243 319
rect 236 315 239 317
rect 241 315 243 317
rect 236 313 243 315
rect 254 314 259 317
rect 236 310 241 313
rect 252 312 259 314
rect 252 310 254 312
rect 256 310 259 312
rect 208 308 211 310
rect 213 308 215 310
rect 208 306 215 308
rect 86 298 88 300
rect 90 298 93 300
rect 86 296 93 298
rect 149 298 152 300
rect 154 298 156 300
rect 149 296 156 298
rect 190 300 197 306
rect 252 308 259 310
rect 261 308 272 317
rect 263 306 272 308
rect 274 306 279 317
rect 281 312 286 317
rect 281 310 288 312
rect 377 311 382 318
rect 281 308 284 310
rect 286 308 288 310
rect 281 306 288 308
rect 375 309 382 311
rect 375 307 377 309
rect 379 307 382 309
rect 190 298 192 300
rect 194 298 197 300
rect 190 296 197 298
rect 263 300 270 306
rect 375 305 382 307
rect 384 305 389 318
rect 391 305 396 318
rect 398 309 409 318
rect 411 316 418 318
rect 411 314 414 316
rect 416 314 418 316
rect 411 312 418 314
rect 428 312 433 317
rect 411 309 416 312
rect 426 310 433 312
rect 398 305 407 309
rect 400 300 407 305
rect 426 308 428 310
rect 430 308 433 310
rect 426 306 433 308
rect 435 306 440 317
rect 442 308 453 317
rect 455 314 460 317
rect 470 314 481 319
rect 455 312 462 314
rect 455 310 458 312
rect 460 310 462 312
rect 470 312 472 314
rect 474 312 481 314
rect 470 310 481 312
rect 483 317 490 319
rect 483 315 486 317
rect 488 315 490 317
rect 483 313 490 315
rect 502 314 507 317
rect 483 310 488 313
rect 500 312 507 314
rect 500 310 502 312
rect 504 310 507 312
rect 455 308 462 310
rect 442 306 451 308
rect 263 298 265 300
rect 267 298 270 300
rect 263 296 270 298
rect 400 298 403 300
rect 405 298 407 300
rect 400 296 407 298
rect 444 300 451 306
rect 500 308 507 310
rect 509 308 520 317
rect 511 306 520 308
rect 522 306 527 317
rect 529 312 534 317
rect 555 312 560 317
rect 529 310 536 312
rect 529 308 532 310
rect 534 308 536 310
rect 529 306 536 308
rect 553 310 560 312
rect 553 308 555 310
rect 557 308 560 310
rect 553 306 560 308
rect 562 306 567 317
rect 569 308 580 317
rect 582 314 587 317
rect 582 312 589 314
rect 604 312 609 317
rect 582 310 585 312
rect 587 310 589 312
rect 582 308 589 310
rect 602 310 609 312
rect 602 308 604 310
rect 606 308 609 310
rect 569 306 578 308
rect 444 298 447 300
rect 449 298 451 300
rect 444 296 451 298
rect 511 300 518 306
rect 511 298 513 300
rect 515 298 518 300
rect 511 296 518 298
rect 571 300 578 306
rect 602 306 609 308
rect 611 306 616 317
rect 618 308 629 317
rect 631 314 636 317
rect 631 312 638 314
rect 631 310 634 312
rect 636 310 638 312
rect 631 308 638 310
rect 645 310 652 312
rect 645 308 647 310
rect 649 308 652 310
rect 618 306 627 308
rect 571 298 574 300
rect 576 298 578 300
rect 571 296 578 298
rect 620 300 627 306
rect 645 306 652 308
rect 620 298 623 300
rect 625 298 627 300
rect 620 296 627 298
rect 647 300 652 306
rect 654 300 659 312
rect 661 304 673 312
rect 661 302 669 304
rect 671 302 673 304
rect 661 300 673 302
rect 85 288 91 290
rect 85 286 87 288
rect 89 286 91 288
rect 85 284 91 286
rect 69 281 74 284
rect 45 279 54 281
rect 45 277 47 279
rect 49 277 54 279
rect 45 276 54 277
rect 33 273 38 276
rect 31 271 38 273
rect 31 269 33 271
rect 35 269 38 271
rect 31 267 38 269
rect 40 272 54 276
rect 56 276 64 281
rect 56 274 59 276
rect 61 274 64 276
rect 56 272 64 274
rect 66 278 74 281
rect 66 276 69 278
rect 71 276 74 278
rect 66 272 74 276
rect 76 272 81 284
rect 83 272 91 284
rect 126 282 131 286
rect 104 279 111 282
rect 104 277 106 279
rect 108 277 111 279
rect 104 275 111 277
rect 40 267 45 272
rect 106 267 111 275
rect 113 271 121 282
rect 113 269 116 271
rect 118 269 121 271
rect 113 267 121 269
rect 123 279 131 282
rect 123 277 126 279
rect 128 277 131 279
rect 123 272 131 277
rect 123 270 126 272
rect 128 270 131 272
rect 123 267 131 270
rect 133 280 140 286
rect 177 288 184 290
rect 177 286 180 288
rect 182 286 184 288
rect 133 278 136 280
rect 138 278 140 280
rect 177 280 184 286
rect 159 278 166 280
rect 133 267 142 278
rect 144 273 149 278
rect 159 276 161 278
rect 163 276 166 278
rect 159 274 166 276
rect 144 271 151 273
rect 144 269 147 271
rect 149 269 151 271
rect 161 269 166 274
rect 168 269 173 280
rect 175 278 184 280
rect 257 288 263 290
rect 257 286 259 288
rect 261 286 263 288
rect 257 284 263 286
rect 461 288 468 290
rect 461 286 463 288
rect 465 286 468 288
rect 241 281 246 284
rect 217 279 226 281
rect 175 269 186 278
rect 188 276 195 278
rect 217 277 219 279
rect 221 277 226 279
rect 217 276 226 277
rect 188 274 191 276
rect 193 274 195 276
rect 188 272 195 274
rect 205 273 210 276
rect 188 269 193 272
rect 203 271 210 273
rect 203 269 205 271
rect 207 269 210 271
rect 144 267 151 269
rect 203 267 210 269
rect 212 272 226 276
rect 228 276 236 281
rect 228 274 231 276
rect 233 274 236 276
rect 228 272 236 274
rect 238 278 246 281
rect 238 276 241 278
rect 243 276 246 278
rect 238 272 246 276
rect 248 272 253 284
rect 255 272 263 284
rect 461 280 468 286
rect 548 288 554 290
rect 548 286 550 288
rect 552 286 554 288
rect 548 284 554 286
rect 592 288 599 290
rect 592 286 595 288
rect 597 286 599 288
rect 532 281 537 284
rect 461 278 470 280
rect 450 276 457 278
rect 273 273 278 276
rect 212 267 217 272
rect 271 271 278 273
rect 271 269 273 271
rect 275 269 278 271
rect 271 267 278 269
rect 280 274 291 276
rect 280 272 287 274
rect 289 272 291 274
rect 450 274 452 276
rect 454 274 457 276
rect 450 272 457 274
rect 280 267 291 272
rect 452 269 457 272
rect 459 269 470 278
rect 472 269 477 280
rect 479 278 486 280
rect 479 276 482 278
rect 484 276 486 278
rect 508 279 517 281
rect 508 277 510 279
rect 512 277 517 279
rect 508 276 517 277
rect 479 274 486 276
rect 479 269 484 274
rect 496 273 501 276
rect 494 271 501 273
rect 494 269 496 271
rect 498 269 501 271
rect 494 267 501 269
rect 503 272 517 276
rect 519 276 527 281
rect 519 274 522 276
rect 524 274 527 276
rect 519 272 527 274
rect 529 278 537 281
rect 529 276 532 278
rect 534 276 537 278
rect 529 272 537 276
rect 539 272 544 284
rect 546 272 554 284
rect 592 280 599 286
rect 668 288 674 290
rect 668 286 670 288
rect 672 286 674 288
rect 574 278 581 280
rect 574 276 576 278
rect 578 276 581 278
rect 574 274 581 276
rect 503 267 508 272
rect 576 269 581 274
rect 583 269 588 280
rect 590 278 599 280
rect 590 269 601 278
rect 603 276 610 278
rect 668 281 674 286
rect 657 279 664 281
rect 657 278 659 279
rect 646 276 653 278
rect 603 274 606 276
rect 608 274 610 276
rect 603 272 610 274
rect 618 274 629 276
rect 618 272 620 274
rect 622 272 629 274
rect 603 269 608 272
rect 618 267 629 272
rect 631 273 636 276
rect 646 274 648 276
rect 650 274 653 276
rect 631 271 638 273
rect 631 269 634 271
rect 636 269 638 271
rect 646 270 653 274
rect 655 277 659 278
rect 661 277 664 279
rect 655 273 664 277
rect 666 280 674 281
rect 666 276 677 280
rect 666 273 674 276
rect 655 270 660 273
rect 631 267 638 269
rect 81 170 92 175
rect 32 159 40 170
rect 32 157 35 159
rect 37 157 40 159
rect 32 155 40 157
rect 42 166 50 170
rect 42 164 45 166
rect 47 164 50 166
rect 42 155 50 164
rect 52 166 60 170
rect 81 168 83 170
rect 85 168 92 170
rect 52 164 55 166
rect 57 164 60 166
rect 52 159 60 164
rect 52 157 55 159
rect 57 157 60 159
rect 52 155 60 157
rect 81 166 92 168
rect 94 173 101 175
rect 94 171 97 173
rect 99 171 101 173
rect 94 169 101 171
rect 113 170 118 173
rect 94 166 99 169
rect 111 168 118 170
rect 111 166 113 168
rect 115 166 118 168
rect 111 164 118 166
rect 120 164 131 173
rect 122 162 131 164
rect 133 162 138 173
rect 140 168 145 173
rect 446 172 453 174
rect 446 170 448 172
rect 450 170 453 172
rect 140 166 147 168
rect 140 164 143 166
rect 145 164 147 166
rect 140 162 147 164
rect 122 156 129 162
rect 156 159 164 170
rect 156 157 159 159
rect 161 157 164 159
rect 122 154 124 156
rect 126 154 129 156
rect 156 155 164 157
rect 166 166 174 170
rect 166 164 169 166
rect 171 164 174 166
rect 166 155 174 164
rect 176 166 184 170
rect 446 168 453 170
rect 176 164 179 166
rect 181 164 184 166
rect 176 159 184 164
rect 176 157 179 159
rect 181 157 184 159
rect 176 155 184 157
rect 448 165 453 168
rect 455 165 466 174
rect 457 161 466 165
rect 468 161 473 174
rect 475 161 480 174
rect 482 167 487 174
rect 482 165 489 167
rect 482 163 485 165
rect 487 163 489 165
rect 482 161 489 163
rect 506 165 513 167
rect 506 163 508 165
rect 510 163 513 165
rect 506 161 513 163
rect 122 152 129 154
rect 457 156 464 161
rect 508 157 513 161
rect 515 157 525 167
rect 527 165 535 167
rect 527 163 530 165
rect 532 163 535 165
rect 527 157 535 163
rect 537 157 546 167
rect 457 154 459 156
rect 461 154 464 156
rect 457 152 464 154
rect 517 156 523 157
rect 517 154 519 156
rect 521 154 523 156
rect 517 152 523 154
rect 539 156 546 157
rect 539 154 541 156
rect 543 154 546 156
rect 539 152 546 154
rect 578 166 587 175
rect 578 164 580 166
rect 582 164 587 166
rect 578 159 587 164
rect 578 157 580 159
rect 582 157 587 159
rect 578 155 587 157
rect 589 155 594 175
rect 596 167 601 175
rect 660 170 665 175
rect 596 165 603 167
rect 596 163 599 165
rect 601 163 603 165
rect 596 161 603 163
rect 596 155 601 161
rect 614 158 622 170
rect 624 158 629 170
rect 631 166 639 170
rect 631 164 634 166
rect 636 164 639 166
rect 631 161 639 164
rect 641 168 649 170
rect 641 166 644 168
rect 646 166 649 168
rect 641 161 649 166
rect 651 166 665 170
rect 667 173 674 175
rect 667 171 670 173
rect 672 171 674 173
rect 667 169 674 171
rect 667 166 672 169
rect 651 165 660 166
rect 651 163 656 165
rect 658 163 660 165
rect 651 161 660 163
rect 631 158 636 161
rect 614 156 620 158
rect 614 154 616 156
rect 618 154 620 156
rect 614 152 620 154
rect 85 144 91 146
rect 85 142 87 144
rect 89 142 91 144
rect 155 144 162 146
rect 85 140 91 142
rect 69 137 74 140
rect 45 135 54 137
rect 45 133 47 135
rect 49 133 54 135
rect 45 132 54 133
rect 33 129 38 132
rect 31 127 38 129
rect 31 125 33 127
rect 35 125 38 127
rect 31 123 38 125
rect 40 128 54 132
rect 56 132 64 137
rect 56 130 59 132
rect 61 130 64 132
rect 56 128 64 130
rect 66 134 74 137
rect 66 132 69 134
rect 71 132 74 134
rect 66 128 74 132
rect 76 128 81 140
rect 83 128 91 140
rect 104 137 109 143
rect 102 135 109 137
rect 102 133 104 135
rect 106 133 109 135
rect 102 131 109 133
rect 40 123 45 128
rect 104 123 109 131
rect 111 123 116 143
rect 118 141 127 143
rect 155 142 158 144
rect 160 142 162 144
rect 118 139 123 141
rect 125 139 127 141
rect 118 134 127 139
rect 155 136 162 142
rect 471 144 477 146
rect 471 142 473 144
rect 475 142 477 144
rect 548 144 555 146
rect 548 142 551 144
rect 553 142 555 144
rect 118 132 123 134
rect 125 132 127 134
rect 118 123 127 132
rect 137 134 144 136
rect 137 132 139 134
rect 141 132 144 134
rect 137 130 144 132
rect 139 125 144 130
rect 146 125 151 136
rect 153 134 162 136
rect 153 125 164 134
rect 166 132 173 134
rect 166 130 169 132
rect 171 130 173 132
rect 166 128 173 130
rect 187 129 192 132
rect 166 125 171 128
rect 185 127 192 129
rect 185 125 187 127
rect 189 125 192 127
rect 185 123 192 125
rect 194 130 205 132
rect 194 128 201 130
rect 203 128 205 130
rect 194 123 205 128
rect 471 137 477 142
rect 548 137 555 142
rect 592 144 599 146
rect 592 142 595 144
rect 597 142 599 144
rect 450 135 457 137
rect 450 133 452 135
rect 454 133 457 135
rect 450 131 457 133
rect 459 135 467 137
rect 459 133 462 135
rect 464 133 467 135
rect 459 131 467 133
rect 469 131 479 137
rect 481 135 489 137
rect 481 133 484 135
rect 486 133 489 135
rect 481 131 489 133
rect 491 135 498 137
rect 491 133 494 135
rect 496 133 498 135
rect 491 131 498 133
rect 523 135 530 137
rect 523 133 525 135
rect 527 133 530 135
rect 523 131 530 133
rect 525 124 530 131
rect 532 124 537 137
rect 539 124 544 137
rect 546 133 555 137
rect 592 136 599 142
rect 646 141 655 143
rect 646 139 648 141
rect 650 139 655 141
rect 574 134 581 136
rect 546 124 557 133
rect 559 130 564 133
rect 574 132 576 134
rect 578 132 581 134
rect 574 130 581 132
rect 559 128 566 130
rect 559 126 562 128
rect 564 126 566 128
rect 559 124 566 126
rect 576 125 581 130
rect 583 125 588 136
rect 590 134 599 136
rect 590 125 601 134
rect 603 132 610 134
rect 646 134 655 139
rect 646 132 648 134
rect 650 132 655 134
rect 603 130 606 132
rect 608 130 610 132
rect 603 128 610 130
rect 618 130 629 132
rect 618 128 620 130
rect 622 128 629 130
rect 603 125 608 128
rect 618 123 629 128
rect 631 129 636 132
rect 631 127 638 129
rect 631 125 634 127
rect 636 125 638 127
rect 631 123 638 125
rect 646 123 655 132
rect 657 123 662 143
rect 664 137 669 143
rect 664 135 671 137
rect 664 133 667 135
rect 669 133 671 135
rect 664 131 671 133
rect 664 123 669 131
rect 79 26 90 31
rect 32 15 40 26
rect 32 13 35 15
rect 37 13 40 15
rect 32 11 40 13
rect 42 22 50 26
rect 42 20 45 22
rect 47 20 50 22
rect 42 11 50 20
rect 52 22 60 26
rect 79 24 81 26
rect 83 24 90 26
rect 52 20 55 22
rect 57 20 60 22
rect 52 15 60 20
rect 52 13 55 15
rect 57 13 60 15
rect 52 11 60 13
rect 79 22 90 24
rect 92 29 99 31
rect 92 27 95 29
rect 97 27 99 29
rect 92 25 99 27
rect 156 26 161 31
rect 92 22 97 25
rect 110 14 118 26
rect 120 14 125 26
rect 127 22 135 26
rect 127 20 130 22
rect 132 20 135 22
rect 127 17 135 20
rect 137 24 145 26
rect 137 22 140 24
rect 142 22 145 24
rect 137 17 145 22
rect 147 22 161 26
rect 163 29 170 31
rect 163 27 166 29
rect 168 27 170 29
rect 163 25 170 27
rect 180 25 188 31
rect 163 22 168 25
rect 180 23 182 25
rect 184 23 188 25
rect 147 21 156 22
rect 147 19 152 21
rect 154 19 156 21
rect 180 21 188 23
rect 190 29 198 31
rect 190 27 193 29
rect 195 27 198 29
rect 190 21 198 27
rect 200 22 208 31
rect 376 26 387 31
rect 376 24 378 26
rect 380 24 387 26
rect 376 22 387 24
rect 389 29 396 31
rect 389 27 392 29
rect 394 27 396 29
rect 389 25 396 27
rect 389 22 394 25
rect 200 21 204 22
rect 147 17 156 19
rect 127 14 132 17
rect 110 12 116 14
rect 110 10 112 12
rect 114 10 116 12
rect 110 8 116 10
rect 202 20 204 21
rect 206 20 208 22
rect 202 18 208 20
rect 411 12 420 31
rect 411 10 414 12
rect 416 11 420 12
rect 422 11 427 31
rect 429 11 434 31
rect 436 11 441 31
rect 443 23 448 31
rect 512 26 517 31
rect 443 21 450 23
rect 443 19 446 21
rect 448 19 450 21
rect 443 17 450 19
rect 443 11 448 17
rect 466 14 474 26
rect 476 14 481 26
rect 483 22 491 26
rect 483 20 486 22
rect 488 20 491 22
rect 483 17 491 20
rect 493 24 501 26
rect 493 22 496 24
rect 498 22 501 24
rect 493 17 501 22
rect 503 22 517 26
rect 519 29 526 31
rect 519 27 522 29
rect 524 27 526 29
rect 519 25 526 27
rect 519 22 524 25
rect 536 24 541 29
rect 534 22 541 24
rect 503 21 512 22
rect 503 19 508 21
rect 510 19 512 21
rect 503 17 512 19
rect 534 20 536 22
rect 538 20 541 22
rect 534 18 541 20
rect 543 18 548 29
rect 550 20 561 29
rect 563 26 568 29
rect 563 24 570 26
rect 563 22 566 24
rect 568 22 570 24
rect 563 20 570 22
rect 578 24 585 28
rect 578 22 580 24
rect 582 22 585 24
rect 578 20 585 22
rect 587 25 592 28
rect 660 26 665 31
rect 587 21 596 25
rect 587 20 591 21
rect 550 18 559 20
rect 483 14 488 17
rect 466 12 472 14
rect 416 10 418 11
rect 411 8 418 10
rect 466 10 468 12
rect 470 10 472 12
rect 466 8 472 10
rect 552 12 559 18
rect 589 19 591 20
rect 593 19 596 21
rect 589 17 596 19
rect 598 17 606 25
rect 552 10 555 12
rect 557 10 559 12
rect 552 8 559 10
rect 600 12 606 17
rect 600 10 602 12
rect 604 10 606 12
rect 600 8 606 10
rect 614 14 622 26
rect 624 14 629 26
rect 631 22 639 26
rect 631 20 634 22
rect 636 20 639 22
rect 631 17 639 20
rect 641 24 649 26
rect 641 22 644 24
rect 646 22 649 24
rect 641 17 649 22
rect 651 22 665 26
rect 667 29 674 31
rect 667 27 670 29
rect 672 27 674 29
rect 667 25 674 27
rect 667 22 672 25
rect 651 21 660 22
rect 651 19 656 21
rect 658 19 660 21
rect 651 17 660 19
rect 631 14 636 17
rect 614 12 620 14
rect 614 10 616 12
rect 618 10 620 12
rect 614 8 620 10
<< pdif >>
rect 39 684 46 686
rect 39 682 41 684
rect 43 682 46 684
rect 39 680 46 682
rect 41 659 46 680
rect 48 670 62 686
rect 48 668 51 670
rect 53 668 62 670
rect 64 684 72 686
rect 64 682 67 684
rect 69 682 72 684
rect 64 677 72 682
rect 64 675 67 677
rect 69 675 72 677
rect 64 668 72 675
rect 74 677 82 686
rect 74 675 77 677
rect 79 675 82 677
rect 74 668 82 675
rect 48 663 60 668
rect 48 661 51 663
rect 53 661 60 663
rect 48 659 60 661
rect 77 659 82 668
rect 84 671 89 686
rect 104 679 109 687
rect 102 677 109 679
rect 102 675 104 677
rect 106 675 109 677
rect 84 669 91 671
rect 84 667 87 669
rect 89 667 91 669
rect 84 665 91 667
rect 102 670 109 675
rect 102 668 104 670
rect 106 668 109 670
rect 102 666 109 668
rect 84 659 89 665
rect 104 659 109 666
rect 111 659 116 687
rect 118 670 127 687
rect 135 684 142 686
rect 135 682 137 684
rect 139 682 142 684
rect 135 677 142 682
rect 135 675 137 677
rect 139 675 142 677
rect 135 673 142 675
rect 118 668 123 670
rect 125 668 127 670
rect 137 668 142 673
rect 144 679 150 686
rect 187 684 194 686
rect 187 682 189 684
rect 191 682 194 684
rect 187 680 194 682
rect 144 672 152 679
rect 144 670 147 672
rect 149 670 152 672
rect 144 668 152 670
rect 118 663 127 668
rect 146 666 152 668
rect 154 677 162 679
rect 154 675 157 677
rect 159 675 162 677
rect 154 670 162 675
rect 154 668 157 670
rect 159 668 162 670
rect 154 666 162 668
rect 164 670 171 679
rect 164 668 167 670
rect 169 668 171 670
rect 164 666 171 668
rect 118 661 123 663
rect 125 661 127 663
rect 118 659 127 661
rect 189 659 194 680
rect 196 670 210 686
rect 196 668 199 670
rect 201 668 210 670
rect 212 684 220 686
rect 212 682 215 684
rect 217 682 220 684
rect 212 677 220 682
rect 212 675 215 677
rect 217 675 220 677
rect 212 668 220 675
rect 222 677 230 686
rect 222 675 225 677
rect 227 675 230 677
rect 222 668 230 675
rect 196 663 208 668
rect 196 661 199 663
rect 201 661 208 663
rect 196 659 208 661
rect 225 659 230 668
rect 232 671 237 686
rect 309 685 316 687
rect 309 683 311 685
rect 313 683 316 685
rect 232 669 239 671
rect 232 667 235 669
rect 237 667 239 669
rect 232 665 239 667
rect 249 667 256 680
rect 249 665 251 667
rect 253 665 256 667
rect 232 659 237 665
rect 249 663 256 665
rect 258 677 266 680
rect 258 675 261 677
rect 263 675 266 677
rect 258 670 266 675
rect 258 668 261 670
rect 263 668 266 670
rect 258 663 266 668
rect 268 667 276 680
rect 268 665 271 667
rect 273 665 276 667
rect 268 663 276 665
rect 278 677 286 680
rect 278 675 281 677
rect 283 675 286 677
rect 278 670 286 675
rect 278 668 281 670
rect 283 668 286 670
rect 278 663 286 668
rect 288 663 296 680
rect 309 678 316 683
rect 309 676 311 678
rect 313 676 316 678
rect 309 674 316 676
rect 311 669 316 674
rect 318 670 327 687
rect 318 669 322 670
rect 320 668 322 669
rect 324 668 327 670
rect 320 666 327 668
rect 497 671 505 684
rect 497 669 500 671
rect 502 669 505 671
rect 497 664 505 669
rect 290 660 296 663
rect 497 662 500 664
rect 502 662 505 664
rect 290 658 292 660
rect 294 658 296 660
rect 290 656 296 658
rect 497 660 505 662
rect 507 678 515 684
rect 507 676 510 678
rect 512 676 515 678
rect 507 668 515 676
rect 517 679 525 684
rect 543 684 550 686
rect 543 682 545 684
rect 547 682 550 684
rect 543 680 550 682
rect 517 677 520 679
rect 522 677 525 679
rect 517 672 525 677
rect 517 670 520 672
rect 522 670 525 672
rect 517 668 525 670
rect 507 660 512 668
rect 545 659 550 680
rect 552 670 566 686
rect 552 668 555 670
rect 557 668 566 670
rect 568 684 576 686
rect 568 682 571 684
rect 573 682 576 684
rect 568 677 576 682
rect 568 675 571 677
rect 573 675 576 677
rect 568 668 576 675
rect 578 677 586 686
rect 578 675 581 677
rect 583 675 586 677
rect 578 668 586 675
rect 552 663 564 668
rect 552 661 555 663
rect 557 661 564 663
rect 552 659 564 661
rect 581 659 586 668
rect 588 671 593 686
rect 606 685 613 687
rect 606 683 608 685
rect 610 683 613 685
rect 606 678 613 683
rect 606 676 608 678
rect 610 676 613 678
rect 606 674 613 676
rect 588 669 595 671
rect 608 669 613 674
rect 615 670 624 687
rect 615 669 619 670
rect 588 667 591 669
rect 593 667 595 669
rect 588 665 595 667
rect 588 659 593 665
rect 617 668 619 669
rect 621 668 624 670
rect 617 666 624 668
rect 634 670 641 686
rect 634 668 636 670
rect 638 668 641 670
rect 634 663 641 668
rect 634 661 636 663
rect 638 661 641 663
rect 634 659 641 661
rect 643 659 648 686
rect 650 684 658 686
rect 650 682 653 684
rect 655 682 658 684
rect 650 677 658 682
rect 650 675 653 677
rect 655 675 658 677
rect 650 659 658 675
rect 660 659 665 686
rect 667 670 674 686
rect 667 668 670 670
rect 672 668 674 670
rect 667 663 674 668
rect 667 661 670 663
rect 672 661 674 663
rect 667 659 674 661
rect 31 645 38 647
rect 31 643 33 645
rect 35 643 38 645
rect 31 638 38 643
rect 31 636 33 638
rect 35 636 38 638
rect 31 623 38 636
rect 40 638 48 647
rect 40 636 43 638
rect 45 636 48 638
rect 40 631 48 636
rect 40 629 43 631
rect 45 629 48 631
rect 40 623 48 629
rect 50 645 58 647
rect 50 643 53 645
rect 55 643 58 645
rect 170 648 176 650
rect 170 646 172 648
rect 174 646 176 648
rect 50 638 58 643
rect 50 636 53 638
rect 55 636 58 638
rect 78 638 85 640
rect 106 638 112 640
rect 78 637 80 638
rect 50 623 58 636
rect 69 632 74 637
rect 67 630 74 632
rect 67 628 69 630
rect 71 628 74 630
rect 67 623 74 628
rect 67 621 69 623
rect 71 621 74 623
rect 67 619 74 621
rect 76 636 80 637
rect 82 636 85 638
rect 76 619 85 636
rect 97 633 102 638
rect 95 631 102 633
rect 95 629 97 631
rect 99 629 102 631
rect 95 624 102 629
rect 95 622 97 624
rect 99 622 102 624
rect 95 620 102 622
rect 104 636 112 638
rect 104 634 107 636
rect 109 634 112 636
rect 104 627 112 634
rect 114 638 122 640
rect 114 636 117 638
rect 119 636 122 638
rect 114 631 122 636
rect 114 629 117 631
rect 119 629 122 631
rect 114 627 122 629
rect 124 638 131 640
rect 170 639 176 646
rect 209 648 216 650
rect 209 646 212 648
rect 214 646 216 648
rect 209 645 216 646
rect 124 636 127 638
rect 129 636 131 638
rect 124 627 131 636
rect 141 634 146 639
rect 139 632 146 634
rect 139 630 141 632
rect 143 630 146 632
rect 104 620 110 627
rect 139 625 146 630
rect 139 623 141 625
rect 143 623 146 625
rect 139 621 146 623
rect 148 637 156 639
rect 148 635 151 637
rect 153 635 156 637
rect 148 626 156 635
rect 158 637 166 639
rect 158 635 161 637
rect 163 635 166 637
rect 158 630 166 635
rect 158 628 161 630
rect 163 628 166 630
rect 158 626 166 628
rect 168 638 176 639
rect 168 626 178 638
rect 148 621 154 626
rect 173 625 178 626
rect 180 636 187 638
rect 180 634 183 636
rect 185 634 187 636
rect 180 629 187 634
rect 180 627 183 629
rect 185 627 187 629
rect 180 625 187 627
rect 209 620 218 645
rect 220 620 225 645
rect 227 620 232 645
rect 234 620 239 645
rect 241 638 246 645
rect 579 645 587 647
rect 502 638 509 640
rect 241 630 249 638
rect 241 628 244 630
rect 246 628 249 630
rect 241 620 249 628
rect 251 620 256 638
rect 258 620 263 638
rect 265 620 270 638
rect 272 636 279 638
rect 272 634 275 636
rect 277 634 279 636
rect 272 629 279 634
rect 272 627 275 629
rect 277 627 279 629
rect 272 620 279 627
rect 502 636 505 638
rect 507 637 509 638
rect 579 643 582 645
rect 584 643 587 645
rect 543 638 549 640
rect 507 636 511 637
rect 502 619 511 636
rect 513 632 518 637
rect 534 633 539 638
rect 513 630 520 632
rect 513 628 516 630
rect 518 628 520 630
rect 513 623 520 628
rect 513 621 516 623
rect 518 621 520 623
rect 513 619 520 621
rect 532 631 539 633
rect 532 629 534 631
rect 536 629 539 631
rect 532 624 539 629
rect 532 622 534 624
rect 536 622 539 624
rect 532 620 539 622
rect 541 636 549 638
rect 541 634 544 636
rect 546 634 549 636
rect 541 627 549 634
rect 551 638 559 640
rect 551 636 554 638
rect 556 636 559 638
rect 551 631 559 636
rect 551 629 554 631
rect 556 629 559 631
rect 551 627 559 629
rect 561 638 568 640
rect 561 636 564 638
rect 566 636 568 638
rect 561 627 568 636
rect 579 638 587 643
rect 579 636 582 638
rect 584 636 587 638
rect 541 620 547 627
rect 579 623 587 636
rect 589 638 597 647
rect 589 636 592 638
rect 594 636 597 638
rect 589 631 597 636
rect 589 629 592 631
rect 594 629 597 631
rect 589 623 597 629
rect 599 645 606 647
rect 599 643 602 645
rect 604 643 606 645
rect 599 638 606 643
rect 616 641 621 647
rect 599 636 602 638
rect 604 636 606 638
rect 599 623 606 636
rect 614 639 621 641
rect 614 637 616 639
rect 618 637 621 639
rect 614 635 621 637
rect 616 620 621 635
rect 623 638 628 647
rect 645 645 657 647
rect 645 643 652 645
rect 654 643 657 645
rect 645 638 657 643
rect 623 631 631 638
rect 623 629 626 631
rect 628 629 631 631
rect 623 620 631 629
rect 633 631 641 638
rect 633 629 636 631
rect 638 629 641 631
rect 633 624 641 629
rect 633 622 636 624
rect 638 622 641 624
rect 633 620 641 622
rect 643 636 652 638
rect 654 636 657 638
rect 643 620 657 636
rect 659 626 664 647
rect 659 624 666 626
rect 659 622 662 624
rect 664 622 666 624
rect 659 620 666 622
rect 39 540 46 542
rect 39 538 41 540
rect 43 538 46 540
rect 39 536 46 538
rect 41 515 46 536
rect 48 526 62 542
rect 48 524 51 526
rect 53 524 62 526
rect 64 540 72 542
rect 64 538 67 540
rect 69 538 72 540
rect 64 533 72 538
rect 64 531 67 533
rect 69 531 72 533
rect 64 524 72 531
rect 74 533 82 542
rect 74 531 77 533
rect 79 531 82 533
rect 74 524 82 531
rect 48 519 60 524
rect 48 517 51 519
rect 53 517 60 519
rect 48 515 60 517
rect 77 515 82 524
rect 84 527 89 542
rect 84 525 91 527
rect 84 523 87 525
rect 89 523 91 525
rect 84 521 91 523
rect 99 526 106 539
rect 99 524 101 526
rect 103 524 106 526
rect 84 515 89 521
rect 99 519 106 524
rect 99 517 101 519
rect 103 517 106 519
rect 99 515 106 517
rect 108 533 116 539
rect 108 531 111 533
rect 113 531 116 533
rect 108 526 116 531
rect 108 524 111 526
rect 113 524 116 526
rect 108 515 116 524
rect 118 526 126 539
rect 118 524 121 526
rect 123 524 126 526
rect 118 519 126 524
rect 118 517 121 519
rect 123 517 126 519
rect 118 515 126 517
rect 143 526 150 543
rect 143 524 145 526
rect 147 524 150 526
rect 143 519 150 524
rect 143 517 145 519
rect 147 517 150 519
rect 143 515 150 517
rect 152 515 157 543
rect 159 515 164 543
rect 166 533 174 543
rect 166 531 169 533
rect 171 531 174 533
rect 166 526 174 531
rect 166 524 169 526
rect 171 524 174 526
rect 166 515 174 524
rect 176 515 181 543
rect 183 515 188 543
rect 190 526 197 543
rect 190 524 193 526
rect 195 524 197 526
rect 211 535 218 537
rect 211 533 213 535
rect 215 533 218 535
rect 211 528 218 533
rect 211 526 213 528
rect 215 526 218 528
rect 211 524 218 526
rect 220 536 225 537
rect 442 541 449 543
rect 244 536 250 541
rect 220 524 230 536
rect 190 519 197 524
rect 222 523 230 524
rect 232 534 240 536
rect 232 532 235 534
rect 237 532 240 534
rect 232 527 240 532
rect 232 525 235 527
rect 237 525 240 527
rect 232 523 240 525
rect 242 527 250 536
rect 242 525 245 527
rect 247 525 250 527
rect 242 523 250 525
rect 252 539 259 541
rect 252 537 255 539
rect 257 537 259 539
rect 252 532 259 537
rect 252 530 255 532
rect 257 530 259 532
rect 442 539 444 541
rect 446 539 449 541
rect 442 534 449 539
rect 442 532 444 534
rect 446 532 449 534
rect 442 530 449 532
rect 252 528 259 530
rect 252 523 257 528
rect 444 525 449 530
rect 451 526 460 543
rect 451 525 455 526
rect 190 517 193 519
rect 195 517 197 519
rect 190 515 197 517
rect 222 516 228 523
rect 453 524 455 525
rect 457 524 460 526
rect 453 522 460 524
rect 510 526 517 542
rect 510 524 512 526
rect 514 524 517 526
rect 510 519 517 524
rect 222 514 224 516
rect 226 514 228 516
rect 222 512 228 514
rect 510 517 512 519
rect 514 517 517 519
rect 510 515 517 517
rect 519 515 524 542
rect 526 540 534 542
rect 526 538 529 540
rect 531 538 534 540
rect 526 533 534 538
rect 526 531 529 533
rect 531 531 534 533
rect 526 515 534 531
rect 536 515 541 542
rect 543 526 550 542
rect 579 535 585 542
rect 543 524 546 526
rect 548 524 550 526
rect 543 519 550 524
rect 558 526 565 535
rect 558 524 560 526
rect 562 524 565 526
rect 558 522 565 524
rect 567 533 575 535
rect 567 531 570 533
rect 572 531 575 533
rect 567 526 575 531
rect 567 524 570 526
rect 572 524 575 526
rect 567 522 575 524
rect 577 528 585 535
rect 577 526 580 528
rect 582 526 585 528
rect 577 524 585 526
rect 587 540 594 542
rect 587 538 590 540
rect 592 538 594 540
rect 587 533 594 538
rect 587 531 590 533
rect 592 531 594 533
rect 587 529 594 531
rect 604 541 611 543
rect 604 539 606 541
rect 608 539 611 541
rect 604 534 611 539
rect 604 532 606 534
rect 608 532 611 534
rect 604 530 611 532
rect 587 524 592 529
rect 606 525 611 530
rect 613 526 622 543
rect 613 525 617 526
rect 577 522 583 524
rect 543 517 546 519
rect 548 517 550 519
rect 615 524 617 525
rect 619 524 622 526
rect 615 522 622 524
rect 634 526 641 542
rect 634 524 636 526
rect 638 524 641 526
rect 634 519 641 524
rect 543 515 550 517
rect 634 517 636 519
rect 638 517 641 519
rect 634 515 641 517
rect 643 515 648 542
rect 650 540 658 542
rect 650 538 653 540
rect 655 538 658 540
rect 650 533 658 538
rect 650 531 653 533
rect 655 531 658 533
rect 650 515 658 531
rect 660 515 665 542
rect 667 526 674 542
rect 667 524 670 526
rect 672 524 674 526
rect 667 519 674 524
rect 667 517 670 519
rect 672 517 674 519
rect 667 515 674 517
rect 36 496 41 503
rect 34 494 41 496
rect 34 492 36 494
rect 38 492 41 494
rect 34 487 41 492
rect 34 485 36 487
rect 38 485 41 487
rect 34 483 41 485
rect 36 475 41 483
rect 43 475 48 503
rect 50 501 59 503
rect 50 499 55 501
rect 57 499 59 501
rect 50 494 59 499
rect 50 492 55 494
rect 57 492 59 494
rect 78 494 85 496
rect 153 497 158 503
rect 106 494 112 496
rect 78 493 80 494
rect 50 475 59 492
rect 69 488 74 493
rect 67 486 74 488
rect 67 484 69 486
rect 71 484 74 486
rect 67 479 74 484
rect 67 477 69 479
rect 71 477 74 479
rect 67 475 74 477
rect 76 492 80 493
rect 82 492 85 494
rect 76 475 85 492
rect 97 489 102 494
rect 95 487 102 489
rect 95 485 97 487
rect 99 485 102 487
rect 95 480 102 485
rect 95 478 97 480
rect 99 478 102 480
rect 95 476 102 478
rect 104 492 112 494
rect 104 490 107 492
rect 109 490 112 492
rect 104 483 112 490
rect 114 494 122 496
rect 114 492 117 494
rect 119 492 122 494
rect 114 487 122 492
rect 114 485 117 487
rect 119 485 122 487
rect 114 483 122 485
rect 124 494 131 496
rect 124 492 127 494
rect 129 492 131 494
rect 124 483 131 492
rect 151 495 158 497
rect 151 493 153 495
rect 155 493 158 495
rect 151 491 158 493
rect 104 476 110 483
rect 153 476 158 491
rect 160 494 165 503
rect 182 501 194 503
rect 182 499 189 501
rect 191 499 194 501
rect 182 494 194 499
rect 160 487 168 494
rect 160 485 163 487
rect 165 485 168 487
rect 160 476 168 485
rect 170 487 178 494
rect 170 485 173 487
rect 175 485 178 487
rect 170 480 178 485
rect 170 478 173 480
rect 175 478 178 480
rect 170 476 178 478
rect 180 492 189 494
rect 191 492 194 494
rect 180 476 194 492
rect 196 482 201 503
rect 219 494 226 496
rect 219 492 221 494
rect 223 492 226 494
rect 219 483 226 492
rect 228 494 236 496
rect 228 492 231 494
rect 233 492 236 494
rect 228 487 236 492
rect 228 485 231 487
rect 233 485 236 487
rect 228 483 236 485
rect 238 494 244 496
rect 444 497 449 503
rect 442 495 449 497
rect 238 492 246 494
rect 238 490 241 492
rect 243 490 246 492
rect 238 483 246 490
rect 196 480 203 482
rect 196 478 199 480
rect 201 478 203 480
rect 196 476 203 478
rect 240 476 246 483
rect 248 489 253 494
rect 442 493 444 495
rect 446 493 449 495
rect 442 491 449 493
rect 248 487 255 489
rect 248 485 251 487
rect 253 485 255 487
rect 248 480 255 485
rect 248 478 251 480
rect 253 478 255 480
rect 248 476 255 478
rect 444 476 449 491
rect 451 494 456 503
rect 473 501 485 503
rect 473 499 480 501
rect 482 499 485 501
rect 473 494 485 499
rect 451 487 459 494
rect 451 485 454 487
rect 456 485 459 487
rect 451 476 459 485
rect 461 487 469 494
rect 461 485 464 487
rect 466 485 469 487
rect 461 480 469 485
rect 461 478 464 480
rect 466 478 469 480
rect 461 476 469 478
rect 471 492 480 494
rect 482 492 485 494
rect 471 476 485 492
rect 487 482 492 503
rect 521 494 527 496
rect 512 489 517 494
rect 510 487 517 489
rect 510 485 512 487
rect 514 485 517 487
rect 487 480 494 482
rect 510 480 517 485
rect 487 478 490 480
rect 492 478 494 480
rect 487 476 494 478
rect 510 478 512 480
rect 514 478 517 480
rect 510 476 517 478
rect 519 492 527 494
rect 519 490 522 492
rect 524 490 527 492
rect 519 483 527 490
rect 529 494 537 496
rect 529 492 532 494
rect 534 492 537 494
rect 529 487 537 492
rect 529 485 532 487
rect 534 485 537 487
rect 529 483 537 485
rect 539 494 546 496
rect 616 497 621 503
rect 614 495 621 497
rect 539 492 542 494
rect 544 492 546 494
rect 539 483 546 492
rect 554 492 562 494
rect 554 490 557 492
rect 559 490 562 492
rect 519 476 525 483
rect 554 476 562 490
rect 564 487 572 494
rect 564 485 567 487
rect 569 485 572 487
rect 564 480 572 485
rect 564 478 567 480
rect 569 478 572 480
rect 564 476 572 478
rect 574 492 582 494
rect 574 490 577 492
rect 579 490 582 492
rect 574 485 582 490
rect 574 483 577 485
rect 579 483 582 485
rect 574 476 582 483
rect 584 487 592 494
rect 584 485 587 487
rect 589 485 592 487
rect 584 480 592 485
rect 584 478 587 480
rect 589 478 592 480
rect 584 476 592 478
rect 594 492 602 494
rect 594 490 597 492
rect 599 490 602 492
rect 614 493 616 495
rect 618 493 621 495
rect 614 491 621 493
rect 594 485 602 490
rect 594 483 597 485
rect 599 483 602 485
rect 594 476 602 483
rect 616 476 621 491
rect 623 494 628 503
rect 645 501 657 503
rect 645 499 652 501
rect 654 499 657 501
rect 645 494 657 499
rect 623 487 631 494
rect 623 485 626 487
rect 628 485 631 487
rect 623 476 631 485
rect 633 487 641 494
rect 633 485 636 487
rect 638 485 641 487
rect 633 480 641 485
rect 633 478 636 480
rect 638 478 641 480
rect 633 476 641 478
rect 643 492 652 494
rect 654 492 657 494
rect 643 476 657 492
rect 659 482 664 503
rect 659 480 666 482
rect 659 478 662 480
rect 664 478 666 480
rect 659 476 666 478
rect 67 396 74 398
rect 67 394 69 396
rect 71 394 74 396
rect 32 391 40 394
rect 32 389 34 391
rect 36 389 40 391
rect 32 384 40 389
rect 32 382 34 384
rect 36 382 40 384
rect 32 380 40 382
rect 42 391 50 394
rect 42 389 45 391
rect 47 389 50 391
rect 42 384 50 389
rect 42 382 45 384
rect 47 382 50 384
rect 42 380 50 382
rect 52 382 60 394
rect 52 380 56 382
rect 58 380 60 382
rect 67 389 74 394
rect 67 387 69 389
rect 71 387 74 389
rect 67 380 74 387
rect 76 391 82 398
rect 116 396 123 398
rect 116 394 118 396
rect 120 394 123 396
rect 76 384 84 391
rect 76 382 79 384
rect 81 382 84 384
rect 76 380 84 382
rect 54 378 60 380
rect 78 378 84 380
rect 86 389 94 391
rect 86 387 89 389
rect 91 387 94 389
rect 86 382 94 387
rect 86 380 89 382
rect 91 380 94 382
rect 86 378 94 380
rect 96 382 103 391
rect 116 389 123 394
rect 116 387 118 389
rect 120 387 123 389
rect 116 385 123 387
rect 96 380 99 382
rect 101 380 103 382
rect 118 380 123 385
rect 125 391 131 398
rect 190 391 196 398
rect 125 384 133 391
rect 125 382 128 384
rect 130 382 133 384
rect 125 380 133 382
rect 96 378 103 380
rect 127 378 133 380
rect 135 389 143 391
rect 135 387 138 389
rect 140 387 143 389
rect 135 382 143 387
rect 135 380 138 382
rect 140 380 143 382
rect 135 378 143 380
rect 145 382 152 391
rect 145 380 148 382
rect 150 380 152 382
rect 145 378 152 380
rect 169 382 176 391
rect 169 380 171 382
rect 173 380 176 382
rect 169 378 176 380
rect 178 389 186 391
rect 178 387 181 389
rect 183 387 186 389
rect 178 382 186 387
rect 178 380 181 382
rect 183 380 186 382
rect 178 378 186 380
rect 188 384 196 391
rect 188 382 191 384
rect 193 382 196 384
rect 188 380 196 382
rect 198 396 205 398
rect 198 394 201 396
rect 203 394 205 396
rect 198 389 205 394
rect 198 387 201 389
rect 203 387 205 389
rect 198 385 205 387
rect 215 397 222 399
rect 215 395 217 397
rect 219 395 222 397
rect 215 390 222 395
rect 215 388 217 390
rect 219 388 222 390
rect 215 386 222 388
rect 198 380 203 385
rect 217 381 222 386
rect 224 382 233 399
rect 243 396 250 398
rect 243 394 245 396
rect 247 394 250 396
rect 243 389 250 394
rect 243 387 245 389
rect 247 387 250 389
rect 243 385 250 387
rect 224 381 228 382
rect 188 378 194 380
rect 226 380 228 381
rect 230 380 233 382
rect 245 380 250 385
rect 252 391 258 398
rect 287 395 294 397
rect 287 393 289 395
rect 291 393 294 395
rect 252 384 260 391
rect 252 382 255 384
rect 257 382 260 384
rect 252 380 260 382
rect 226 378 233 380
rect 254 378 260 380
rect 262 389 270 391
rect 262 387 265 389
rect 267 387 270 389
rect 262 382 270 387
rect 262 380 265 382
rect 267 380 270 382
rect 262 378 270 380
rect 272 382 279 391
rect 287 388 294 393
rect 287 386 289 388
rect 291 386 294 388
rect 287 384 294 386
rect 272 380 275 382
rect 277 380 279 382
rect 272 378 279 380
rect 289 379 294 384
rect 296 392 302 397
rect 321 392 326 393
rect 296 383 304 392
rect 296 381 299 383
rect 301 381 304 383
rect 296 379 304 381
rect 306 390 314 392
rect 306 388 309 390
rect 311 388 314 390
rect 306 383 314 388
rect 306 381 309 383
rect 311 381 314 383
rect 306 379 314 381
rect 316 380 326 392
rect 328 391 335 393
rect 438 391 444 398
rect 328 389 331 391
rect 333 389 335 391
rect 328 384 335 389
rect 328 382 331 384
rect 333 382 335 384
rect 328 380 335 382
rect 417 382 424 391
rect 417 380 419 382
rect 421 380 424 382
rect 316 379 324 380
rect 318 372 324 379
rect 417 378 424 380
rect 426 389 434 391
rect 426 387 429 389
rect 431 387 434 389
rect 426 382 434 387
rect 426 380 429 382
rect 431 380 434 382
rect 426 378 434 380
rect 436 384 444 391
rect 436 382 439 384
rect 441 382 444 384
rect 436 380 444 382
rect 446 396 453 398
rect 446 394 449 396
rect 451 394 453 396
rect 446 389 453 394
rect 446 387 449 389
rect 451 387 453 389
rect 446 385 453 387
rect 462 397 469 399
rect 462 395 464 397
rect 466 395 469 397
rect 462 390 469 395
rect 462 388 464 390
rect 466 388 469 390
rect 462 386 469 388
rect 446 380 451 385
rect 464 381 469 386
rect 471 382 480 399
rect 511 391 517 398
rect 471 381 475 382
rect 436 378 442 380
rect 318 370 320 372
rect 322 370 324 372
rect 318 368 324 370
rect 473 380 475 381
rect 477 380 480 382
rect 473 378 480 380
rect 490 382 497 391
rect 490 380 492 382
rect 494 380 497 382
rect 490 378 497 380
rect 499 389 507 391
rect 499 387 502 389
rect 504 387 507 389
rect 499 382 507 387
rect 499 380 502 382
rect 504 380 507 382
rect 499 378 507 380
rect 509 384 517 391
rect 509 382 512 384
rect 514 382 517 384
rect 509 380 517 382
rect 519 396 526 398
rect 519 394 522 396
rect 524 394 526 396
rect 519 389 526 394
rect 519 387 522 389
rect 524 387 526 389
rect 519 385 526 387
rect 538 396 545 398
rect 538 394 540 396
rect 542 394 545 396
rect 538 389 545 394
rect 538 387 540 389
rect 542 387 545 389
rect 538 385 545 387
rect 519 380 524 385
rect 540 380 545 385
rect 547 391 553 398
rect 582 391 589 393
rect 547 384 555 391
rect 547 382 550 384
rect 552 382 555 384
rect 547 380 555 382
rect 509 378 515 380
rect 549 378 555 380
rect 557 389 565 391
rect 557 387 560 389
rect 562 387 565 389
rect 557 382 565 387
rect 557 380 560 382
rect 562 380 565 382
rect 557 378 565 380
rect 567 382 574 391
rect 567 380 570 382
rect 572 380 574 382
rect 582 389 584 391
rect 586 389 589 391
rect 582 384 589 389
rect 582 382 584 384
rect 586 382 589 384
rect 582 380 589 382
rect 591 392 596 393
rect 615 392 621 397
rect 591 380 601 392
rect 567 378 574 380
rect 593 379 601 380
rect 603 390 611 392
rect 603 388 606 390
rect 608 388 611 390
rect 603 383 611 388
rect 603 381 606 383
rect 608 381 611 383
rect 603 379 611 381
rect 613 383 621 392
rect 613 381 616 383
rect 618 381 621 383
rect 613 379 621 381
rect 623 395 630 397
rect 623 393 626 395
rect 628 393 630 395
rect 623 388 630 393
rect 623 386 626 388
rect 628 386 630 388
rect 623 384 630 386
rect 623 379 628 384
rect 638 382 645 391
rect 638 380 640 382
rect 642 380 645 382
rect 593 372 599 379
rect 638 375 645 380
rect 593 370 595 372
rect 597 370 599 372
rect 638 373 640 375
rect 642 373 645 375
rect 638 371 645 373
rect 647 389 655 391
rect 647 387 650 389
rect 652 387 655 389
rect 647 382 655 387
rect 647 380 650 382
rect 652 380 655 382
rect 647 371 655 380
rect 657 382 665 391
rect 657 380 660 382
rect 662 380 665 382
rect 657 375 665 380
rect 657 373 660 375
rect 662 373 665 375
rect 657 371 665 373
rect 667 389 674 391
rect 667 387 670 389
rect 672 387 674 389
rect 667 382 674 387
rect 667 380 670 382
rect 672 380 674 382
rect 667 378 674 380
rect 667 371 672 378
rect 593 368 599 370
rect 106 360 112 362
rect 33 352 38 359
rect 31 350 38 352
rect 31 348 33 350
rect 35 348 38 350
rect 31 343 38 348
rect 31 341 33 343
rect 35 341 38 343
rect 31 339 38 341
rect 40 357 48 359
rect 40 355 43 357
rect 45 355 48 357
rect 40 350 48 355
rect 40 348 43 350
rect 45 348 48 350
rect 40 339 48 348
rect 50 350 58 359
rect 50 348 53 350
rect 55 348 58 350
rect 50 343 58 348
rect 50 341 53 343
rect 55 341 58 343
rect 50 339 58 341
rect 60 357 67 359
rect 60 355 63 357
rect 65 355 67 357
rect 106 358 108 360
rect 110 358 112 360
rect 60 350 67 355
rect 106 351 112 358
rect 60 348 63 350
rect 65 348 67 350
rect 60 339 67 348
rect 77 346 82 351
rect 75 344 82 346
rect 75 342 77 344
rect 79 342 82 344
rect 75 337 82 342
rect 75 335 77 337
rect 79 335 82 337
rect 75 333 82 335
rect 84 349 92 351
rect 84 347 87 349
rect 89 347 92 349
rect 84 338 92 347
rect 94 349 102 351
rect 94 347 97 349
rect 99 347 102 349
rect 94 342 102 347
rect 94 340 97 342
rect 99 340 102 342
rect 94 338 102 340
rect 104 350 112 351
rect 131 350 138 352
rect 104 338 114 350
rect 84 333 90 338
rect 109 337 114 338
rect 116 348 123 350
rect 116 346 119 348
rect 121 346 123 348
rect 116 341 123 346
rect 116 339 119 341
rect 121 339 123 341
rect 131 348 133 350
rect 135 348 138 350
rect 131 339 138 348
rect 140 350 148 352
rect 140 348 143 350
rect 145 348 148 350
rect 140 343 148 348
rect 140 341 143 343
rect 145 341 148 343
rect 140 339 148 341
rect 150 350 156 352
rect 190 350 196 352
rect 150 348 158 350
rect 150 346 153 348
rect 155 346 158 348
rect 150 339 158 346
rect 116 337 123 339
rect 152 332 158 339
rect 160 345 165 350
rect 181 345 186 350
rect 160 343 167 345
rect 160 341 163 343
rect 165 341 167 343
rect 160 336 167 341
rect 160 334 163 336
rect 165 334 167 336
rect 160 332 167 334
rect 179 343 186 345
rect 179 341 181 343
rect 183 341 186 343
rect 179 336 186 341
rect 179 334 181 336
rect 183 334 186 336
rect 179 332 186 334
rect 188 348 196 350
rect 188 346 191 348
rect 193 346 196 348
rect 188 339 196 346
rect 198 350 206 352
rect 198 348 201 350
rect 203 348 206 350
rect 198 343 206 348
rect 198 341 201 343
rect 203 341 206 343
rect 198 339 206 341
rect 208 350 215 352
rect 208 348 211 350
rect 213 348 215 350
rect 208 339 215 348
rect 225 350 232 352
rect 225 348 228 350
rect 230 349 232 350
rect 381 360 387 362
rect 381 358 383 360
rect 385 358 387 360
rect 263 350 269 352
rect 230 348 234 349
rect 188 332 194 339
rect 225 331 234 348
rect 236 344 241 349
rect 254 345 259 350
rect 236 342 243 344
rect 236 340 239 342
rect 241 340 243 342
rect 236 335 243 340
rect 236 333 239 335
rect 241 333 243 335
rect 236 331 243 333
rect 252 343 259 345
rect 252 341 254 343
rect 256 341 259 343
rect 252 336 259 341
rect 252 334 254 336
rect 256 334 259 336
rect 252 332 259 334
rect 261 348 269 350
rect 261 346 264 348
rect 266 346 269 348
rect 261 339 269 346
rect 271 350 279 352
rect 271 348 274 350
rect 276 348 279 350
rect 271 343 279 348
rect 271 341 274 343
rect 276 341 279 343
rect 271 339 279 341
rect 281 350 288 352
rect 381 351 387 358
rect 381 350 389 351
rect 281 348 284 350
rect 286 348 288 350
rect 281 339 288 348
rect 370 348 377 350
rect 370 346 372 348
rect 374 346 377 348
rect 370 341 377 346
rect 370 339 372 341
rect 374 339 377 341
rect 261 332 267 339
rect 370 337 377 339
rect 379 338 389 350
rect 391 349 399 351
rect 391 347 394 349
rect 396 347 399 349
rect 391 342 399 347
rect 391 340 394 342
rect 396 340 399 342
rect 391 338 399 340
rect 401 349 409 351
rect 401 347 404 349
rect 406 347 409 349
rect 401 338 409 347
rect 379 337 384 338
rect 403 333 409 338
rect 411 346 416 351
rect 426 350 433 352
rect 426 348 428 350
rect 430 348 433 350
rect 411 344 418 346
rect 411 342 414 344
rect 416 342 418 344
rect 411 337 418 342
rect 426 339 433 348
rect 435 350 443 352
rect 435 348 438 350
rect 440 348 443 350
rect 435 343 443 348
rect 435 341 438 343
rect 440 341 443 343
rect 435 339 443 341
rect 445 350 451 352
rect 472 350 479 352
rect 445 348 453 350
rect 445 346 448 348
rect 450 346 453 348
rect 445 339 453 346
rect 411 335 414 337
rect 416 335 418 337
rect 411 333 418 335
rect 447 332 453 339
rect 455 345 460 350
rect 472 348 475 350
rect 477 349 479 350
rect 511 350 517 352
rect 477 348 481 349
rect 455 343 462 345
rect 455 341 458 343
rect 460 341 462 343
rect 455 336 462 341
rect 455 334 458 336
rect 460 334 462 336
rect 455 332 462 334
rect 472 331 481 348
rect 483 344 488 349
rect 502 345 507 350
rect 483 342 490 344
rect 483 340 486 342
rect 488 340 490 342
rect 483 335 490 340
rect 483 333 486 335
rect 488 333 490 335
rect 483 331 490 333
rect 500 343 507 345
rect 500 341 502 343
rect 504 341 507 343
rect 500 336 507 341
rect 500 334 502 336
rect 504 334 507 336
rect 500 332 507 334
rect 509 348 517 350
rect 509 346 512 348
rect 514 346 517 348
rect 509 339 517 346
rect 519 350 527 352
rect 519 348 522 350
rect 524 348 527 350
rect 519 343 527 348
rect 519 341 522 343
rect 524 341 527 343
rect 519 339 527 341
rect 529 350 536 352
rect 529 348 532 350
rect 534 348 536 350
rect 529 339 536 348
rect 553 350 560 352
rect 553 348 555 350
rect 557 348 560 350
rect 553 339 560 348
rect 562 350 570 352
rect 562 348 565 350
rect 567 348 570 350
rect 562 343 570 348
rect 562 341 565 343
rect 567 341 570 343
rect 562 339 570 341
rect 572 350 578 352
rect 602 350 609 352
rect 572 348 580 350
rect 572 346 575 348
rect 577 346 580 348
rect 572 339 580 346
rect 509 332 515 339
rect 574 332 580 339
rect 582 345 587 350
rect 602 348 604 350
rect 606 348 609 350
rect 582 343 589 345
rect 582 341 585 343
rect 587 341 589 343
rect 582 336 589 341
rect 602 339 609 348
rect 611 350 619 352
rect 611 348 614 350
rect 616 348 619 350
rect 611 343 619 348
rect 611 341 614 343
rect 616 341 619 343
rect 611 339 619 341
rect 621 350 627 352
rect 645 350 651 352
rect 621 348 629 350
rect 621 346 624 348
rect 626 346 629 348
rect 621 339 629 346
rect 582 334 585 336
rect 587 334 589 336
rect 582 332 589 334
rect 623 332 629 339
rect 631 343 638 350
rect 631 341 634 343
rect 636 341 638 343
rect 631 336 638 341
rect 645 348 647 350
rect 649 348 653 350
rect 645 336 653 348
rect 655 348 663 350
rect 655 346 658 348
rect 660 346 663 348
rect 655 341 663 346
rect 655 339 658 341
rect 660 339 663 341
rect 655 336 663 339
rect 665 348 673 350
rect 665 346 669 348
rect 671 346 673 348
rect 665 341 673 346
rect 665 339 669 341
rect 671 339 673 341
rect 665 336 673 339
rect 631 334 634 336
rect 636 334 638 336
rect 631 332 638 334
rect 39 252 46 254
rect 39 250 41 252
rect 43 250 46 252
rect 39 248 46 250
rect 41 227 46 248
rect 48 238 62 254
rect 48 236 51 238
rect 53 236 62 238
rect 64 252 72 254
rect 64 250 67 252
rect 69 250 72 252
rect 64 245 72 250
rect 64 243 67 245
rect 69 243 72 245
rect 64 236 72 243
rect 74 245 82 254
rect 74 243 77 245
rect 79 243 82 245
rect 74 236 82 243
rect 48 231 60 236
rect 48 229 51 231
rect 53 229 60 231
rect 48 227 60 229
rect 77 227 82 236
rect 84 239 89 254
rect 103 247 111 254
rect 103 245 106 247
rect 108 245 111 247
rect 103 240 111 245
rect 84 237 91 239
rect 84 235 87 237
rect 89 235 91 237
rect 103 238 106 240
rect 108 238 111 240
rect 103 236 111 238
rect 113 252 121 254
rect 113 250 116 252
rect 118 250 121 252
rect 113 245 121 250
rect 113 243 116 245
rect 118 243 121 245
rect 113 236 121 243
rect 123 247 131 254
rect 123 245 126 247
rect 128 245 131 247
rect 123 240 131 245
rect 123 238 126 240
rect 128 238 131 240
rect 123 236 131 238
rect 133 252 141 254
rect 133 250 136 252
rect 138 250 141 252
rect 133 245 141 250
rect 133 243 136 245
rect 138 243 141 245
rect 133 236 141 243
rect 143 240 151 254
rect 180 247 186 254
rect 143 238 146 240
rect 148 238 151 240
rect 143 236 151 238
rect 159 238 166 247
rect 159 236 161 238
rect 163 236 166 238
rect 84 233 91 235
rect 84 227 89 233
rect 159 234 166 236
rect 168 245 176 247
rect 168 243 171 245
rect 173 243 176 245
rect 168 238 176 243
rect 168 236 171 238
rect 173 236 176 238
rect 168 234 176 236
rect 178 240 186 247
rect 178 238 181 240
rect 183 238 186 240
rect 178 236 186 238
rect 188 252 195 254
rect 188 250 191 252
rect 193 250 195 252
rect 211 252 218 254
rect 211 250 213 252
rect 215 250 218 252
rect 188 245 195 250
rect 211 248 218 250
rect 188 243 191 245
rect 193 243 195 245
rect 188 241 195 243
rect 188 236 193 241
rect 178 234 184 236
rect 213 227 218 248
rect 220 238 234 254
rect 220 236 223 238
rect 225 236 234 238
rect 236 252 244 254
rect 236 250 239 252
rect 241 250 244 252
rect 236 245 244 250
rect 236 243 239 245
rect 241 243 244 245
rect 236 236 244 243
rect 246 245 254 254
rect 246 243 249 245
rect 251 243 254 245
rect 246 236 254 243
rect 220 231 232 236
rect 220 229 223 231
rect 225 229 232 231
rect 220 227 232 229
rect 249 227 254 236
rect 256 239 261 254
rect 271 253 278 255
rect 271 251 273 253
rect 275 251 278 253
rect 271 246 278 251
rect 271 244 273 246
rect 275 244 278 246
rect 271 242 278 244
rect 256 237 263 239
rect 273 237 278 242
rect 280 238 289 255
rect 450 252 457 254
rect 450 250 452 252
rect 454 250 457 252
rect 450 245 457 250
rect 450 243 452 245
rect 454 243 457 245
rect 450 241 457 243
rect 280 237 284 238
rect 256 235 259 237
rect 261 235 263 237
rect 256 233 263 235
rect 256 227 261 233
rect 282 236 284 237
rect 286 236 289 238
rect 452 236 457 241
rect 459 247 465 254
rect 502 252 509 254
rect 502 250 504 252
rect 506 250 509 252
rect 502 248 509 250
rect 459 240 467 247
rect 459 238 462 240
rect 464 238 467 240
rect 459 236 467 238
rect 282 234 289 236
rect 461 234 467 236
rect 469 245 477 247
rect 469 243 472 245
rect 474 243 477 245
rect 469 238 477 243
rect 469 236 472 238
rect 474 236 477 238
rect 469 234 477 236
rect 479 238 486 247
rect 479 236 482 238
rect 484 236 486 238
rect 479 234 486 236
rect 504 227 509 248
rect 511 238 525 254
rect 511 236 514 238
rect 516 236 525 238
rect 527 252 535 254
rect 527 250 530 252
rect 532 250 535 252
rect 527 245 535 250
rect 527 243 530 245
rect 532 243 535 245
rect 527 236 535 243
rect 537 245 545 254
rect 537 243 540 245
rect 542 243 545 245
rect 537 236 545 243
rect 511 231 523 236
rect 511 229 514 231
rect 516 229 523 231
rect 511 227 523 229
rect 540 227 545 236
rect 547 239 552 254
rect 595 247 601 254
rect 547 237 554 239
rect 547 235 550 237
rect 552 235 554 237
rect 547 233 554 235
rect 574 238 581 247
rect 574 236 576 238
rect 578 236 581 238
rect 574 234 581 236
rect 583 245 591 247
rect 583 243 586 245
rect 588 243 591 245
rect 583 238 591 243
rect 583 236 586 238
rect 588 236 591 238
rect 583 234 591 236
rect 593 240 601 247
rect 593 238 596 240
rect 598 238 601 240
rect 593 236 601 238
rect 603 252 610 254
rect 603 250 606 252
rect 608 250 610 252
rect 603 245 610 250
rect 603 243 606 245
rect 608 243 610 245
rect 603 241 610 243
rect 603 236 608 241
rect 620 238 629 255
rect 620 236 623 238
rect 625 237 629 238
rect 631 253 638 255
rect 631 251 634 253
rect 636 251 638 253
rect 631 246 638 251
rect 631 244 634 246
rect 636 244 638 246
rect 631 242 638 244
rect 631 237 636 242
rect 646 238 655 255
rect 625 236 627 237
rect 593 234 599 236
rect 547 227 552 233
rect 620 234 627 236
rect 646 236 648 238
rect 650 236 655 238
rect 646 231 655 236
rect 646 229 648 231
rect 650 229 655 231
rect 646 227 655 229
rect 657 227 662 255
rect 664 247 669 255
rect 664 245 671 247
rect 664 243 667 245
rect 669 243 671 245
rect 664 238 671 243
rect 664 236 667 238
rect 669 236 671 238
rect 664 234 671 236
rect 664 227 669 234
rect 31 213 38 215
rect 31 211 33 213
rect 35 211 38 213
rect 31 206 38 211
rect 31 204 33 206
rect 35 204 38 206
rect 31 188 38 204
rect 40 188 45 215
rect 47 199 55 215
rect 47 197 50 199
rect 52 197 55 199
rect 47 192 55 197
rect 47 190 50 192
rect 52 190 55 192
rect 47 188 55 190
rect 57 188 62 215
rect 64 213 71 215
rect 64 211 67 213
rect 69 211 71 213
rect 477 216 483 218
rect 155 213 162 215
rect 64 206 71 211
rect 64 204 67 206
rect 69 204 71 206
rect 64 188 71 204
rect 83 206 90 208
rect 83 204 86 206
rect 88 205 90 206
rect 155 211 157 213
rect 159 211 162 213
rect 122 206 128 208
rect 88 204 92 205
rect 83 187 92 204
rect 94 200 99 205
rect 113 201 118 206
rect 94 198 101 200
rect 94 196 97 198
rect 99 196 101 198
rect 94 191 101 196
rect 94 189 97 191
rect 99 189 101 191
rect 94 187 101 189
rect 111 199 118 201
rect 111 197 113 199
rect 115 197 118 199
rect 111 192 118 197
rect 111 190 113 192
rect 115 190 118 192
rect 111 188 118 190
rect 120 204 128 206
rect 120 202 123 204
rect 125 202 128 204
rect 120 195 128 202
rect 130 206 138 208
rect 130 204 133 206
rect 135 204 138 206
rect 130 199 138 204
rect 130 197 133 199
rect 135 197 138 199
rect 130 195 138 197
rect 140 206 147 208
rect 140 204 143 206
rect 145 204 147 206
rect 140 195 147 204
rect 155 206 162 211
rect 155 204 157 206
rect 159 204 162 206
rect 120 188 126 195
rect 155 188 162 204
rect 164 188 169 215
rect 171 199 179 215
rect 171 197 174 199
rect 176 197 179 199
rect 171 192 179 197
rect 171 190 174 192
rect 176 190 179 192
rect 171 188 179 190
rect 181 188 186 215
rect 188 213 195 215
rect 188 211 191 213
rect 193 211 195 213
rect 477 214 479 216
rect 481 214 483 216
rect 188 206 195 211
rect 477 207 483 214
rect 508 213 515 215
rect 508 211 510 213
rect 512 211 515 213
rect 188 204 191 206
rect 193 204 195 206
rect 188 188 195 204
rect 448 202 453 207
rect 446 200 453 202
rect 446 198 448 200
rect 450 198 453 200
rect 446 193 453 198
rect 446 191 448 193
rect 450 191 453 193
rect 446 189 453 191
rect 455 205 463 207
rect 455 203 458 205
rect 460 203 463 205
rect 455 194 463 203
rect 465 205 473 207
rect 465 203 468 205
rect 470 203 473 205
rect 465 198 473 203
rect 465 196 468 198
rect 470 196 473 198
rect 465 194 473 196
rect 475 206 483 207
rect 508 206 515 211
rect 475 194 485 206
rect 455 189 461 194
rect 480 193 485 194
rect 487 204 494 206
rect 487 202 490 204
rect 492 202 494 204
rect 487 197 494 202
rect 487 195 490 197
rect 492 195 494 197
rect 487 193 494 195
rect 508 204 510 206
rect 512 204 515 206
rect 508 187 515 204
rect 517 187 522 215
rect 524 187 529 215
rect 531 206 539 215
rect 531 204 534 206
rect 536 204 539 206
rect 531 199 539 204
rect 531 197 534 199
rect 536 197 539 199
rect 531 187 539 197
rect 541 187 546 215
rect 548 187 553 215
rect 555 213 562 215
rect 555 211 558 213
rect 560 211 562 213
rect 555 206 562 211
rect 555 204 558 206
rect 560 204 562 206
rect 555 187 562 204
rect 579 213 587 215
rect 579 211 582 213
rect 584 211 587 213
rect 579 206 587 211
rect 579 204 582 206
rect 584 204 587 206
rect 579 191 587 204
rect 589 206 597 215
rect 589 204 592 206
rect 594 204 597 206
rect 589 199 597 204
rect 589 197 592 199
rect 594 197 597 199
rect 589 191 597 197
rect 599 213 606 215
rect 599 211 602 213
rect 604 211 606 213
rect 599 206 606 211
rect 616 209 621 215
rect 599 204 602 206
rect 604 204 606 206
rect 599 191 606 204
rect 614 207 621 209
rect 614 205 616 207
rect 618 205 621 207
rect 614 203 621 205
rect 616 188 621 203
rect 623 206 628 215
rect 645 213 657 215
rect 645 211 652 213
rect 654 211 657 213
rect 645 206 657 211
rect 623 199 631 206
rect 623 197 626 199
rect 628 197 631 199
rect 623 188 631 197
rect 633 199 641 206
rect 633 197 636 199
rect 638 197 641 199
rect 633 192 641 197
rect 633 190 636 192
rect 638 190 641 192
rect 633 188 641 190
rect 643 204 652 206
rect 654 204 657 206
rect 643 188 657 204
rect 659 194 664 215
rect 659 192 666 194
rect 659 190 662 192
rect 664 190 666 192
rect 659 188 666 190
rect 39 108 46 110
rect 39 106 41 108
rect 43 106 46 108
rect 39 104 46 106
rect 41 83 46 104
rect 48 94 62 110
rect 48 92 51 94
rect 53 92 62 94
rect 64 108 72 110
rect 64 106 67 108
rect 69 106 72 108
rect 64 101 72 106
rect 64 99 67 101
rect 69 99 72 101
rect 64 92 72 99
rect 74 101 82 110
rect 74 99 77 101
rect 79 99 82 101
rect 74 92 82 99
rect 48 87 60 92
rect 48 85 51 87
rect 53 85 60 87
rect 48 83 60 85
rect 77 83 82 92
rect 84 95 89 110
rect 84 93 91 95
rect 84 91 87 93
rect 89 91 91 93
rect 84 89 91 91
rect 99 94 106 107
rect 99 92 101 94
rect 103 92 106 94
rect 84 83 89 89
rect 99 87 106 92
rect 99 85 101 87
rect 103 85 106 87
rect 99 83 106 85
rect 108 101 116 107
rect 108 99 111 101
rect 113 99 116 101
rect 108 94 116 99
rect 108 92 111 94
rect 113 92 116 94
rect 108 83 116 92
rect 118 94 126 107
rect 158 103 164 110
rect 118 92 121 94
rect 123 92 126 94
rect 118 87 126 92
rect 137 94 144 103
rect 137 92 139 94
rect 141 92 144 94
rect 137 90 144 92
rect 146 101 154 103
rect 146 99 149 101
rect 151 99 154 101
rect 146 94 154 99
rect 146 92 149 94
rect 151 92 154 94
rect 146 90 154 92
rect 156 96 164 103
rect 156 94 159 96
rect 161 94 164 96
rect 156 92 164 94
rect 166 108 173 110
rect 166 106 169 108
rect 171 106 173 108
rect 166 101 173 106
rect 166 99 169 101
rect 171 99 173 101
rect 166 97 173 99
rect 185 109 192 111
rect 185 107 187 109
rect 189 107 192 109
rect 185 102 192 107
rect 185 100 187 102
rect 189 100 192 102
rect 185 98 192 100
rect 166 92 171 97
rect 187 93 192 98
rect 194 94 203 111
rect 194 93 198 94
rect 156 90 162 92
rect 118 85 121 87
rect 123 85 126 87
rect 196 92 198 93
rect 200 92 203 94
rect 426 103 433 110
rect 426 101 428 103
rect 430 101 433 103
rect 426 96 433 101
rect 426 94 428 96
rect 430 94 433 96
rect 426 92 433 94
rect 435 92 440 110
rect 442 92 447 110
rect 449 92 454 110
rect 456 102 464 110
rect 456 100 459 102
rect 461 100 464 102
rect 456 92 464 100
rect 196 90 203 92
rect 118 83 126 85
rect 459 85 464 92
rect 466 85 471 110
rect 473 85 478 110
rect 480 85 485 110
rect 487 85 496 110
rect 518 103 525 105
rect 518 101 520 103
rect 522 101 525 103
rect 518 96 525 101
rect 518 94 520 96
rect 522 94 525 96
rect 518 92 525 94
rect 527 104 532 105
rect 551 104 557 109
rect 527 92 537 104
rect 529 91 537 92
rect 539 102 547 104
rect 539 100 542 102
rect 544 100 547 102
rect 539 95 547 100
rect 539 93 542 95
rect 544 93 547 95
rect 539 91 547 93
rect 549 95 557 104
rect 549 93 552 95
rect 554 93 557 95
rect 549 91 557 93
rect 559 107 566 109
rect 559 105 562 107
rect 564 105 566 107
rect 559 100 566 105
rect 595 103 601 110
rect 559 98 562 100
rect 564 98 566 100
rect 559 96 566 98
rect 559 91 564 96
rect 574 94 581 103
rect 574 92 576 94
rect 578 92 581 94
rect 489 84 496 85
rect 489 82 491 84
rect 493 82 496 84
rect 489 80 496 82
rect 529 84 535 91
rect 574 90 581 92
rect 583 101 591 103
rect 583 99 586 101
rect 588 99 591 101
rect 583 94 591 99
rect 583 92 586 94
rect 588 92 591 94
rect 583 90 591 92
rect 593 96 601 103
rect 593 94 596 96
rect 598 94 601 96
rect 593 92 601 94
rect 603 108 610 110
rect 603 106 606 108
rect 608 106 610 108
rect 603 101 610 106
rect 603 99 606 101
rect 608 99 610 101
rect 603 97 610 99
rect 603 92 608 97
rect 620 94 629 111
rect 620 92 623 94
rect 625 93 629 94
rect 631 109 638 111
rect 631 107 634 109
rect 636 107 638 109
rect 631 102 638 107
rect 631 100 634 102
rect 636 100 638 102
rect 631 98 638 100
rect 631 93 636 98
rect 647 94 655 107
rect 625 92 627 93
rect 593 90 599 92
rect 620 90 627 92
rect 647 92 650 94
rect 652 92 655 94
rect 647 87 655 92
rect 529 82 531 84
rect 533 82 535 84
rect 529 80 535 82
rect 647 85 650 87
rect 652 85 655 87
rect 647 83 655 85
rect 657 101 665 107
rect 657 99 660 101
rect 662 99 665 101
rect 657 94 665 99
rect 657 92 660 94
rect 662 92 665 94
rect 657 83 665 92
rect 667 94 674 107
rect 667 92 670 94
rect 672 92 674 94
rect 667 87 674 92
rect 667 85 670 87
rect 672 85 674 87
rect 667 83 674 85
rect 31 69 38 71
rect 31 67 33 69
rect 35 67 38 69
rect 31 62 38 67
rect 31 60 33 62
rect 35 60 38 62
rect 31 44 38 60
rect 40 44 45 71
rect 47 55 55 71
rect 47 53 50 55
rect 52 53 55 55
rect 47 48 55 53
rect 47 46 50 48
rect 52 46 55 48
rect 47 44 55 46
rect 57 44 62 71
rect 64 69 71 71
rect 64 67 67 69
rect 69 67 71 69
rect 64 62 71 67
rect 64 60 67 62
rect 69 60 71 62
rect 64 44 71 60
rect 81 62 88 64
rect 81 60 84 62
rect 86 61 88 62
rect 112 65 117 71
rect 110 63 117 65
rect 110 61 112 63
rect 114 61 117 63
rect 86 60 90 61
rect 81 43 90 60
rect 92 56 97 61
rect 110 59 117 61
rect 92 54 99 56
rect 92 52 95 54
rect 97 52 99 54
rect 92 47 99 52
rect 92 45 95 47
rect 97 45 99 47
rect 92 43 99 45
rect 112 44 117 59
rect 119 62 124 71
rect 141 69 153 71
rect 141 67 148 69
rect 150 67 153 69
rect 141 62 153 67
rect 119 55 127 62
rect 119 53 122 55
rect 124 53 127 55
rect 119 44 127 53
rect 129 55 137 62
rect 129 53 132 55
rect 134 53 137 55
rect 129 48 137 53
rect 129 46 132 48
rect 134 46 137 48
rect 129 44 137 46
rect 139 60 148 62
rect 150 60 153 62
rect 139 44 153 60
rect 155 50 160 71
rect 193 62 198 70
rect 180 60 188 62
rect 180 58 183 60
rect 185 58 188 60
rect 180 53 188 58
rect 180 51 183 53
rect 185 51 188 53
rect 155 48 162 50
rect 155 46 158 48
rect 160 46 162 48
rect 155 44 162 46
rect 180 46 188 51
rect 190 54 198 62
rect 190 52 193 54
rect 195 52 198 54
rect 190 46 198 52
rect 200 68 208 70
rect 409 72 415 74
rect 409 70 411 72
rect 413 70 415 72
rect 200 66 203 68
rect 205 66 208 68
rect 409 67 415 70
rect 200 61 208 66
rect 200 59 203 61
rect 205 59 208 61
rect 200 46 208 59
rect 378 62 385 64
rect 378 60 381 62
rect 383 61 385 62
rect 383 60 387 61
rect 378 43 387 60
rect 389 56 394 61
rect 389 54 396 56
rect 389 52 392 54
rect 394 52 396 54
rect 389 47 396 52
rect 409 50 417 67
rect 419 62 427 67
rect 419 60 422 62
rect 424 60 427 62
rect 419 55 427 60
rect 419 53 422 55
rect 424 53 427 55
rect 419 50 427 53
rect 429 65 437 67
rect 429 63 432 65
rect 434 63 437 65
rect 429 50 437 63
rect 439 62 447 67
rect 439 60 442 62
rect 444 60 447 62
rect 439 55 447 60
rect 439 53 442 55
rect 444 53 447 55
rect 439 50 447 53
rect 449 65 456 67
rect 468 65 473 71
rect 449 63 452 65
rect 454 63 456 65
rect 449 50 456 63
rect 466 63 473 65
rect 466 61 468 63
rect 470 61 473 63
rect 466 59 473 61
rect 389 45 392 47
rect 394 45 396 47
rect 389 43 396 45
rect 468 44 473 59
rect 475 62 480 71
rect 497 69 509 71
rect 497 67 504 69
rect 506 67 509 69
rect 497 62 509 67
rect 475 55 483 62
rect 475 53 478 55
rect 480 53 483 55
rect 475 44 483 53
rect 485 55 493 62
rect 485 53 488 55
rect 490 53 493 55
rect 485 48 493 53
rect 485 46 488 48
rect 490 46 493 48
rect 485 44 493 46
rect 495 60 504 62
rect 506 60 509 62
rect 495 44 509 60
rect 511 50 516 71
rect 578 69 587 71
rect 578 67 580 69
rect 582 67 587 69
rect 534 62 541 64
rect 534 60 536 62
rect 538 60 541 62
rect 534 51 541 60
rect 543 62 551 64
rect 543 60 546 62
rect 548 60 551 62
rect 543 55 551 60
rect 543 53 546 55
rect 548 53 551 55
rect 543 51 551 53
rect 553 62 559 64
rect 578 62 587 67
rect 553 60 561 62
rect 553 58 556 60
rect 558 58 561 60
rect 553 51 561 58
rect 511 48 518 50
rect 511 46 514 48
rect 516 46 518 48
rect 511 44 518 46
rect 555 44 561 51
rect 563 57 568 62
rect 578 60 580 62
rect 582 60 587 62
rect 563 55 570 57
rect 563 53 566 55
rect 568 53 570 55
rect 563 48 570 53
rect 563 46 566 48
rect 568 46 570 48
rect 563 44 570 46
rect 578 43 587 60
rect 589 43 594 71
rect 596 64 601 71
rect 616 65 621 71
rect 596 62 603 64
rect 596 60 599 62
rect 601 60 603 62
rect 596 55 603 60
rect 614 63 621 65
rect 614 61 616 63
rect 618 61 621 63
rect 614 59 621 61
rect 596 53 599 55
rect 601 53 603 55
rect 596 51 603 53
rect 596 43 601 51
rect 616 44 621 59
rect 623 62 628 71
rect 645 69 657 71
rect 645 67 652 69
rect 654 67 657 69
rect 645 62 657 67
rect 623 55 631 62
rect 623 53 626 55
rect 628 53 631 55
rect 623 44 631 53
rect 633 55 641 62
rect 633 53 636 55
rect 638 53 641 55
rect 633 48 641 53
rect 633 46 636 48
rect 638 46 641 48
rect 633 44 641 46
rect 643 60 652 62
rect 654 60 657 62
rect 643 44 657 60
rect 659 50 664 71
rect 659 48 666 50
rect 659 46 662 48
rect 664 46 666 48
rect 659 44 666 46
<< alu1 >>
rect 27 720 336 725
rect 27 718 34 720
rect 36 718 87 720
rect 89 718 101 720
rect 103 718 122 720
rect 124 718 138 720
rect 140 718 148 720
rect 150 718 182 720
rect 184 718 235 720
rect 237 718 289 720
rect 291 718 312 720
rect 314 718 324 720
rect 326 718 336 720
rect 27 717 336 718
rect 494 720 678 725
rect 494 718 500 720
rect 502 718 520 720
rect 522 718 538 720
rect 540 718 591 720
rect 593 718 609 720
rect 611 718 621 720
rect 623 718 633 720
rect 635 718 678 720
rect 494 717 678 718
rect 99 711 116 712
rect 67 710 91 711
rect 67 708 69 710
rect 71 708 91 710
rect 67 707 91 708
rect 39 702 52 704
rect 39 700 40 702
rect 42 700 52 702
rect 39 699 52 700
rect 87 703 91 707
rect 39 698 49 699
rect 47 697 49 698
rect 51 697 52 699
rect 31 686 36 688
rect 31 684 33 686
rect 35 684 36 686
rect 31 672 36 684
rect 47 690 52 697
rect 87 701 88 703
rect 90 701 91 703
rect 31 666 43 672
rect 87 679 91 701
rect 75 678 91 679
rect 75 677 84 678
rect 75 675 77 677
rect 79 676 84 677
rect 86 676 91 678
rect 79 675 91 676
rect 75 674 91 675
rect 99 709 112 711
rect 114 709 116 711
rect 99 708 116 709
rect 99 706 111 708
rect 99 678 103 706
rect 135 709 147 712
rect 249 711 261 712
rect 135 708 144 709
rect 135 706 137 708
rect 139 707 144 708
rect 146 707 147 709
rect 139 706 147 707
rect 215 710 239 711
rect 115 703 119 704
rect 115 701 116 703
rect 118 701 119 703
rect 115 698 119 701
rect 115 697 127 698
rect 107 694 111 696
rect 115 695 118 697
rect 120 695 127 697
rect 115 694 127 695
rect 107 692 108 694
rect 110 692 111 694
rect 107 690 111 692
rect 123 690 127 694
rect 107 686 119 690
rect 115 684 116 686
rect 118 684 119 686
rect 115 682 119 684
rect 135 686 139 706
rect 215 708 217 710
rect 219 708 239 710
rect 215 707 239 708
rect 159 700 164 704
rect 159 698 161 700
rect 163 698 164 700
rect 159 695 164 698
rect 135 684 140 686
rect 135 682 137 684
rect 139 682 140 684
rect 99 677 108 678
rect 99 675 104 677
rect 106 675 108 677
rect 99 674 108 675
rect 102 673 108 674
rect 135 677 140 682
rect 135 675 137 677
rect 139 675 140 677
rect 150 694 164 695
rect 150 692 154 694
rect 156 692 164 694
rect 150 691 164 692
rect 187 703 200 704
rect 187 701 188 703
rect 190 701 200 703
rect 187 699 200 701
rect 187 698 197 699
rect 195 697 197 698
rect 199 697 200 699
rect 158 686 171 687
rect 158 684 164 686
rect 166 684 171 686
rect 158 683 171 684
rect 135 673 140 675
rect 102 671 105 673
rect 107 671 108 673
rect 102 670 108 671
rect 102 668 104 670
rect 106 668 108 670
rect 102 667 108 668
rect 167 677 171 683
rect 167 675 168 677
rect 170 675 171 677
rect 167 674 171 675
rect 179 686 184 688
rect 179 684 181 686
rect 183 684 184 686
rect 179 672 184 684
rect 195 690 200 697
rect 179 669 191 672
rect 179 667 186 669
rect 188 667 191 669
rect 179 666 191 667
rect 235 679 239 707
rect 223 677 239 679
rect 223 675 225 677
rect 227 675 239 677
rect 223 674 239 675
rect 249 709 250 711
rect 252 709 257 711
rect 259 709 261 711
rect 249 708 261 709
rect 249 680 253 708
rect 265 704 269 712
rect 257 700 269 704
rect 273 703 277 712
rect 281 706 293 712
rect 273 701 274 703
rect 276 701 277 703
rect 257 697 261 700
rect 257 695 258 697
rect 260 695 261 697
rect 273 696 277 701
rect 289 700 293 706
rect 289 698 290 700
rect 292 698 293 700
rect 257 694 261 695
rect 257 692 258 694
rect 260 692 261 694
rect 257 690 261 692
rect 265 692 277 696
rect 265 687 271 692
rect 265 685 268 687
rect 270 685 271 687
rect 265 682 271 685
rect 281 686 285 696
rect 289 694 293 698
rect 289 692 290 694
rect 292 692 293 694
rect 289 690 293 692
rect 309 703 313 712
rect 571 710 595 711
rect 309 701 311 703
rect 281 685 293 686
rect 281 683 290 685
rect 292 683 293 685
rect 281 682 293 683
rect 249 678 261 680
rect 249 677 285 678
rect 249 675 261 677
rect 263 675 281 677
rect 283 675 285 677
rect 249 674 285 675
rect 280 670 285 674
rect 280 668 281 670
rect 283 668 285 670
rect 280 666 285 668
rect 289 666 293 682
rect 309 685 313 701
rect 571 708 573 710
rect 575 708 595 710
rect 571 707 595 708
rect 317 696 321 704
rect 497 703 517 704
rect 497 701 510 703
rect 512 701 517 703
rect 497 698 517 701
rect 317 695 329 696
rect 317 694 325 695
rect 317 692 318 694
rect 320 693 325 694
rect 327 693 329 695
rect 320 692 329 693
rect 317 690 329 692
rect 309 683 311 685
rect 309 680 313 683
rect 309 678 321 680
rect 309 676 311 678
rect 313 677 321 678
rect 313 676 318 677
rect 309 675 318 676
rect 320 675 321 677
rect 497 679 501 698
rect 521 693 525 696
rect 523 691 525 693
rect 543 699 556 704
rect 543 698 553 699
rect 551 697 553 698
rect 555 697 556 699
rect 521 687 525 691
rect 512 686 525 687
rect 512 684 522 686
rect 524 684 525 686
rect 512 683 525 684
rect 535 686 540 688
rect 535 684 537 686
rect 539 684 540 686
rect 497 678 514 679
rect 497 676 505 678
rect 507 676 510 678
rect 512 676 514 678
rect 497 675 514 676
rect 309 674 321 675
rect 535 672 540 684
rect 551 693 556 697
rect 551 691 552 693
rect 554 691 556 693
rect 551 690 556 691
rect 535 669 547 672
rect 535 667 536 669
rect 538 667 547 669
rect 535 666 547 667
rect 591 679 595 707
rect 579 677 595 679
rect 579 675 581 677
rect 583 675 595 677
rect 579 674 595 675
rect 606 703 610 712
rect 606 701 608 703
rect 606 685 610 701
rect 614 703 618 704
rect 614 701 615 703
rect 617 701 618 703
rect 637 703 642 712
rect 656 710 674 711
rect 656 708 658 710
rect 660 708 661 710
rect 663 708 674 710
rect 656 707 674 708
rect 637 702 664 703
rect 614 696 618 701
rect 637 700 639 702
rect 641 700 661 702
rect 663 700 664 702
rect 637 699 664 700
rect 660 697 661 699
rect 663 697 664 699
rect 614 694 626 696
rect 660 695 664 697
rect 614 692 615 694
rect 617 692 626 694
rect 614 690 626 692
rect 637 694 654 695
rect 637 692 650 694
rect 652 692 654 694
rect 637 691 654 692
rect 606 683 608 685
rect 606 680 610 683
rect 637 685 642 691
rect 670 687 674 707
rect 637 683 638 685
rect 640 683 642 685
rect 637 682 642 683
rect 652 686 674 687
rect 652 684 671 686
rect 673 684 674 686
rect 652 682 653 684
rect 655 683 674 684
rect 655 682 658 683
rect 606 679 618 680
rect 606 678 613 679
rect 606 676 608 678
rect 610 677 613 678
rect 615 677 618 679
rect 610 676 618 677
rect 606 674 618 676
rect 652 677 658 682
rect 652 675 653 677
rect 655 675 658 677
rect 652 673 658 675
rect 27 660 336 661
rect 27 658 67 660
rect 69 658 138 660
rect 140 658 215 660
rect 217 658 292 660
rect 294 658 312 660
rect 314 658 324 660
rect 326 658 336 660
rect 27 653 336 658
rect 494 660 678 661
rect 494 658 519 660
rect 521 658 571 660
rect 573 658 609 660
rect 611 658 621 660
rect 623 658 678 660
rect 27 648 287 653
rect 27 646 70 648
rect 72 646 82 648
rect 84 646 98 648
rect 100 646 172 648
rect 174 646 186 648
rect 188 646 212 648
rect 214 646 252 648
rect 254 646 274 648
rect 276 646 287 648
rect 27 645 287 646
rect 494 648 678 658
rect 494 646 503 648
rect 505 646 515 648
rect 517 646 535 648
rect 537 646 636 648
rect 638 646 678 648
rect 494 645 678 646
rect 31 626 43 632
rect 67 630 79 632
rect 67 628 69 630
rect 71 628 79 630
rect 67 626 79 628
rect 95 631 100 633
rect 95 629 97 631
rect 99 629 100 631
rect 139 632 144 640
rect 95 628 100 629
rect 95 626 96 628
rect 98 626 100 628
rect 31 607 35 626
rect 47 623 59 624
rect 47 621 56 623
rect 58 621 59 623
rect 47 618 59 621
rect 31 605 32 607
rect 34 605 35 607
rect 31 598 35 605
rect 39 614 43 616
rect 57 616 59 618
rect 39 612 40 614
rect 42 612 43 614
rect 39 608 43 612
rect 55 610 59 616
rect 67 623 71 626
rect 67 621 69 623
rect 39 605 51 608
rect 39 603 48 605
rect 50 603 51 605
rect 39 602 51 603
rect 67 605 71 621
rect 95 624 100 626
rect 95 622 97 624
rect 99 622 100 624
rect 95 620 100 622
rect 75 615 87 616
rect 75 614 84 615
rect 75 612 76 614
rect 78 613 84 614
rect 86 613 87 615
rect 78 612 87 613
rect 75 610 87 612
rect 67 603 69 605
rect 31 597 40 598
rect 31 595 36 597
rect 38 595 40 597
rect 31 594 40 595
rect 67 597 71 603
rect 75 602 79 610
rect 67 595 68 597
rect 70 595 71 597
rect 67 594 71 595
rect 95 600 99 620
rect 127 623 131 632
rect 118 622 131 623
rect 118 620 119 622
rect 121 620 124 622
rect 126 620 131 622
rect 118 619 131 620
rect 139 630 141 632
rect 143 631 144 632
rect 143 630 152 631
rect 139 628 149 630
rect 151 628 152 630
rect 139 627 152 628
rect 139 625 143 627
rect 139 623 141 625
rect 110 614 124 615
rect 110 612 114 614
rect 116 612 124 614
rect 110 611 124 612
rect 119 608 124 611
rect 95 598 97 600
rect 99 598 107 600
rect 95 594 107 598
rect 119 606 120 608
rect 122 606 124 608
rect 119 602 124 606
rect 139 604 143 623
rect 170 623 176 631
rect 207 638 267 639
rect 207 636 208 638
rect 210 636 267 638
rect 207 635 267 636
rect 162 622 184 623
rect 162 621 172 622
rect 162 619 168 621
rect 170 620 172 621
rect 174 620 184 622
rect 170 619 184 620
rect 207 615 211 635
rect 215 630 248 631
rect 215 628 216 630
rect 218 628 244 630
rect 246 628 248 630
rect 215 627 248 628
rect 154 614 167 615
rect 154 612 158 614
rect 160 612 167 614
rect 154 611 167 612
rect 139 602 141 604
rect 139 594 143 602
rect 163 605 167 611
rect 178 614 184 615
rect 178 612 180 614
rect 182 612 184 614
rect 178 608 184 612
rect 207 613 209 615
rect 207 611 211 613
rect 163 603 164 605
rect 166 603 167 605
rect 163 602 167 603
rect 171 605 184 608
rect 171 603 181 605
rect 183 603 184 605
rect 171 602 184 603
rect 215 599 219 627
rect 263 623 267 635
rect 508 630 520 632
rect 508 628 513 630
rect 515 628 516 630
rect 518 628 520 630
rect 508 626 520 628
rect 223 622 258 623
rect 223 620 224 622
rect 226 620 258 622
rect 223 619 258 620
rect 263 619 278 623
rect 516 623 520 626
rect 518 621 520 623
rect 223 608 227 619
rect 254 615 258 619
rect 272 615 278 619
rect 223 606 224 608
rect 226 606 227 608
rect 238 607 244 615
rect 254 611 267 615
rect 272 613 274 615
rect 276 613 278 615
rect 272 612 278 613
rect 500 614 512 616
rect 500 613 509 614
rect 263 609 267 611
rect 500 611 505 613
rect 507 612 509 613
rect 511 612 512 614
rect 507 611 512 612
rect 500 610 512 611
rect 263 607 264 609
rect 266 607 267 609
rect 223 604 227 606
rect 233 606 258 607
rect 233 604 235 606
rect 237 604 249 606
rect 251 604 254 606
rect 256 604 258 606
rect 263 605 267 607
rect 271 607 275 608
rect 271 605 272 607
rect 274 605 275 607
rect 233 603 258 604
rect 271 600 275 605
rect 215 597 245 599
rect 215 595 219 597
rect 221 595 241 597
rect 243 595 245 597
rect 215 594 245 595
rect 263 598 275 600
rect 263 596 264 598
rect 266 596 275 598
rect 263 594 275 596
rect 508 602 512 610
rect 516 605 520 621
rect 518 603 520 605
rect 516 594 520 603
rect 532 631 537 633
rect 532 629 534 631
rect 536 629 537 631
rect 532 624 537 629
rect 532 622 534 624
rect 536 622 537 624
rect 532 620 537 622
rect 564 631 568 632
rect 564 629 565 631
rect 567 629 568 631
rect 532 618 533 620
rect 535 618 536 620
rect 532 600 536 618
rect 564 623 568 629
rect 594 626 606 632
rect 555 622 568 623
rect 555 620 561 622
rect 563 620 568 622
rect 555 619 568 620
rect 578 623 590 624
rect 578 621 586 623
rect 588 621 590 623
rect 578 618 590 621
rect 578 616 580 618
rect 547 614 561 615
rect 547 612 551 614
rect 553 612 561 614
rect 547 611 561 612
rect 532 598 534 600
rect 536 598 544 600
rect 532 594 544 598
rect 556 605 561 611
rect 578 610 582 616
rect 594 614 598 616
rect 594 612 595 614
rect 597 612 598 614
rect 594 608 598 612
rect 556 603 558 605
rect 560 603 561 605
rect 556 602 561 603
rect 586 606 598 608
rect 586 604 595 606
rect 597 604 598 606
rect 586 602 598 604
rect 602 598 606 626
rect 597 597 606 598
rect 597 595 599 597
rect 601 595 603 597
rect 605 595 606 597
rect 614 631 630 632
rect 614 629 622 631
rect 624 629 626 631
rect 628 629 630 631
rect 614 627 630 629
rect 614 606 618 627
rect 662 634 674 640
rect 614 604 615 606
rect 617 604 618 606
rect 614 599 618 604
rect 653 609 658 616
rect 669 622 674 634
rect 669 620 670 622
rect 672 620 674 622
rect 669 618 674 620
rect 653 607 654 609
rect 656 608 658 609
rect 656 607 666 608
rect 653 605 666 607
rect 653 603 663 605
rect 665 603 666 605
rect 653 602 666 603
rect 614 598 638 599
rect 614 596 634 598
rect 636 596 638 598
rect 614 595 638 596
rect 597 594 606 595
rect 27 588 287 589
rect 27 586 70 588
rect 72 586 82 588
rect 84 586 98 588
rect 100 586 108 588
rect 110 586 142 588
rect 144 586 152 588
rect 154 586 230 588
rect 232 586 274 588
rect 276 586 287 588
rect 27 581 287 586
rect 494 588 678 589
rect 494 586 503 588
rect 505 586 515 588
rect 517 586 535 588
rect 537 586 545 588
rect 547 586 616 588
rect 618 586 669 588
rect 671 586 678 588
rect 494 581 678 586
rect 27 576 259 581
rect 27 574 34 576
rect 36 574 87 576
rect 89 574 146 576
rect 148 574 162 576
rect 164 574 184 576
rect 186 574 244 576
rect 246 574 254 576
rect 256 574 259 576
rect 27 573 259 574
rect 438 576 678 581
rect 438 574 445 576
rect 447 574 457 576
rect 459 574 509 576
rect 511 574 579 576
rect 581 574 589 576
rect 591 574 607 576
rect 609 574 619 576
rect 621 574 633 576
rect 635 574 678 576
rect 438 573 678 574
rect 99 567 108 568
rect 67 566 91 567
rect 67 564 69 566
rect 71 564 91 566
rect 67 563 91 564
rect 39 558 52 560
rect 39 556 40 558
rect 42 556 52 558
rect 39 555 52 556
rect 39 554 49 555
rect 47 553 49 554
rect 51 553 52 555
rect 31 542 36 544
rect 31 540 33 542
rect 35 540 36 542
rect 31 528 36 540
rect 47 546 52 553
rect 87 557 91 563
rect 87 555 88 557
rect 90 555 91 557
rect 31 522 43 528
rect 87 535 91 555
rect 75 533 91 535
rect 75 531 77 533
rect 79 531 91 533
rect 75 530 91 531
rect 99 565 104 567
rect 106 565 108 567
rect 99 564 108 565
rect 99 536 103 564
rect 154 566 167 568
rect 154 564 155 566
rect 157 564 167 566
rect 171 567 199 568
rect 171 565 173 567
rect 175 565 195 567
rect 197 565 199 567
rect 171 564 199 565
rect 154 563 167 564
rect 107 557 119 560
rect 162 559 167 563
rect 107 555 112 557
rect 114 555 119 557
rect 146 558 158 559
rect 146 556 147 558
rect 149 556 158 558
rect 146 555 155 556
rect 107 554 119 555
rect 154 554 155 555
rect 157 554 158 556
rect 162 558 170 559
rect 162 556 166 558
rect 168 556 170 558
rect 162 555 170 556
rect 177 558 183 560
rect 177 556 178 558
rect 180 556 183 558
rect 107 550 111 554
rect 107 548 108 550
rect 110 548 111 550
rect 107 546 111 548
rect 123 546 127 552
rect 154 551 158 554
rect 177 551 183 556
rect 143 550 150 551
rect 143 548 145 550
rect 147 548 150 550
rect 143 547 150 548
rect 154 547 183 551
rect 187 558 191 560
rect 187 556 188 558
rect 190 556 191 558
rect 125 544 127 546
rect 115 541 127 544
rect 115 539 119 541
rect 121 539 127 541
rect 146 543 150 547
rect 187 543 191 556
rect 146 542 191 543
rect 146 540 188 542
rect 190 540 191 542
rect 146 539 191 540
rect 115 538 127 539
rect 99 533 111 536
rect 195 535 199 564
rect 255 566 259 568
rect 255 564 256 566
rect 258 564 259 566
rect 214 558 227 560
rect 214 556 224 558
rect 226 556 227 558
rect 214 554 227 556
rect 214 550 220 554
rect 214 548 216 550
rect 218 548 220 550
rect 214 547 220 548
rect 231 551 235 560
rect 255 560 259 564
rect 257 558 259 560
rect 231 550 244 551
rect 231 548 238 550
rect 240 548 241 550
rect 243 548 244 550
rect 231 547 244 548
rect 214 541 228 543
rect 230 541 236 543
rect 214 539 236 541
rect 99 531 100 533
rect 102 531 111 533
rect 162 534 199 535
rect 162 533 196 534
rect 162 531 169 533
rect 171 532 196 533
rect 198 532 199 534
rect 171 531 199 532
rect 99 530 111 531
rect 222 534 228 539
rect 222 532 223 534
rect 225 532 228 534
rect 222 531 228 532
rect 255 539 259 558
rect 257 537 259 539
rect 255 535 259 537
rect 246 532 259 535
rect 246 531 255 532
rect 254 530 255 531
rect 257 530 259 532
rect 442 567 446 568
rect 442 565 443 567
rect 445 565 446 567
rect 442 559 446 565
rect 442 557 444 559
rect 442 541 446 557
rect 450 552 454 560
rect 513 559 518 568
rect 532 566 550 567
rect 532 564 534 566
rect 536 564 550 566
rect 532 563 550 564
rect 513 558 540 559
rect 513 556 515 558
rect 517 556 537 558
rect 539 556 540 558
rect 513 555 540 556
rect 536 553 537 555
rect 539 553 540 555
rect 450 551 462 552
rect 536 551 540 553
rect 450 550 459 551
rect 450 548 451 550
rect 453 549 459 550
rect 461 549 462 551
rect 453 548 462 549
rect 450 546 462 548
rect 486 550 530 551
rect 486 548 487 550
rect 489 548 526 550
rect 528 548 530 550
rect 486 547 530 548
rect 442 539 444 541
rect 442 536 446 539
rect 513 538 518 547
rect 546 543 550 563
rect 565 558 570 560
rect 565 556 567 558
rect 569 556 570 558
rect 565 551 570 556
rect 582 564 594 568
rect 582 562 590 564
rect 592 562 594 564
rect 565 550 579 551
rect 565 548 573 550
rect 575 548 579 550
rect 565 547 579 548
rect 528 540 550 543
rect 528 538 529 540
rect 531 539 550 540
rect 558 542 571 543
rect 558 540 559 542
rect 561 540 563 542
rect 565 540 571 542
rect 558 539 571 540
rect 531 538 534 539
rect 528 536 534 538
rect 442 534 454 536
rect 442 532 444 534
rect 446 532 454 534
rect 442 530 454 532
rect 528 534 529 536
rect 531 534 534 536
rect 528 533 534 534
rect 528 531 529 533
rect 531 531 534 533
rect 254 522 259 530
rect 528 529 534 531
rect 558 530 562 539
rect 590 542 594 562
rect 589 540 594 542
rect 589 538 590 540
rect 592 538 594 540
rect 589 535 594 538
rect 604 559 608 568
rect 604 557 606 559
rect 604 541 608 557
rect 612 552 616 560
rect 637 559 642 568
rect 656 566 674 567
rect 656 564 658 566
rect 660 564 674 566
rect 656 563 674 564
rect 637 558 664 559
rect 637 556 639 558
rect 641 556 646 558
rect 648 556 664 558
rect 637 555 664 556
rect 660 553 661 555
rect 663 553 664 555
rect 612 550 624 552
rect 660 551 664 553
rect 612 548 613 550
rect 615 548 619 550
rect 621 548 624 550
rect 612 546 624 548
rect 637 550 654 551
rect 637 548 650 550
rect 652 548 654 550
rect 637 547 654 548
rect 604 539 606 541
rect 604 538 608 539
rect 604 536 605 538
rect 607 536 608 538
rect 637 541 642 547
rect 670 543 674 563
rect 637 539 638 541
rect 640 539 642 541
rect 637 538 642 539
rect 652 540 674 543
rect 652 538 653 540
rect 655 539 674 540
rect 655 538 658 539
rect 652 537 658 538
rect 589 534 597 535
rect 589 533 594 534
rect 589 531 590 533
rect 592 532 594 533
rect 596 532 597 534
rect 592 531 597 532
rect 604 534 616 536
rect 604 532 606 534
rect 608 532 616 534
rect 589 529 594 531
rect 604 530 616 532
rect 652 535 655 537
rect 657 535 658 537
rect 652 533 658 535
rect 652 531 653 533
rect 655 531 658 533
rect 652 529 658 531
rect 27 516 259 517
rect 27 514 67 516
rect 69 514 210 516
rect 212 514 224 516
rect 226 514 259 516
rect 27 504 259 514
rect 27 502 70 504
rect 72 502 82 504
rect 84 502 98 504
rect 100 502 173 504
rect 175 502 250 504
rect 252 502 259 504
rect 27 501 259 502
rect 438 516 678 517
rect 438 514 445 516
rect 447 514 457 516
rect 459 514 589 516
rect 591 514 607 516
rect 609 514 619 516
rect 621 514 678 516
rect 438 504 678 514
rect 438 502 464 504
rect 466 502 513 504
rect 515 502 557 504
rect 559 502 565 504
rect 567 502 636 504
rect 638 502 678 504
rect 438 501 678 502
rect 34 494 40 495
rect 34 492 36 494
rect 38 492 40 494
rect 34 488 40 492
rect 31 487 40 488
rect 31 485 36 487
rect 38 485 40 487
rect 31 484 40 485
rect 67 486 79 488
rect 67 484 69 486
rect 71 484 79 486
rect 31 461 35 484
rect 67 482 79 484
rect 95 487 100 489
rect 95 485 97 487
rect 99 485 100 487
rect 47 479 59 480
rect 47 477 56 479
rect 58 477 59 479
rect 47 476 59 477
rect 67 479 71 482
rect 67 477 69 479
rect 39 472 51 476
rect 39 470 43 472
rect 39 468 40 470
rect 42 468 43 470
rect 55 471 59 472
rect 55 469 56 471
rect 58 469 59 471
rect 55 468 59 469
rect 39 466 43 468
rect 47 467 59 468
rect 31 459 32 461
rect 34 459 35 461
rect 31 456 35 459
rect 47 465 50 467
rect 52 465 59 467
rect 47 464 59 465
rect 47 458 51 464
rect 67 461 71 477
rect 95 480 100 485
rect 95 478 97 480
rect 99 478 100 480
rect 95 476 100 478
rect 127 486 131 488
rect 127 484 128 486
rect 130 484 131 486
rect 75 470 87 472
rect 75 468 76 470
rect 78 468 87 470
rect 75 466 87 468
rect 67 459 69 461
rect 31 454 43 456
rect 28 453 50 454
rect 28 451 29 453
rect 31 451 44 453
rect 46 451 50 453
rect 28 450 50 451
rect 67 453 71 459
rect 75 461 79 466
rect 75 459 76 461
rect 78 459 79 461
rect 95 462 99 476
rect 95 460 96 462
rect 98 460 99 462
rect 75 458 79 459
rect 67 451 68 453
rect 70 451 71 453
rect 67 450 71 451
rect 95 456 99 460
rect 127 479 131 484
rect 118 478 131 479
rect 118 476 124 478
rect 126 476 131 478
rect 118 475 131 476
rect 151 487 167 488
rect 151 485 163 487
rect 165 485 167 487
rect 151 483 167 485
rect 110 470 124 471
rect 110 468 114 470
rect 116 468 124 470
rect 110 467 124 468
rect 119 463 124 467
rect 95 454 97 456
rect 99 454 107 456
rect 95 450 107 454
rect 119 458 140 463
rect 135 453 140 458
rect 135 451 136 453
rect 138 451 140 453
rect 151 455 155 483
rect 199 494 211 496
rect 199 492 200 494
rect 202 492 211 494
rect 199 490 211 492
rect 190 465 195 472
rect 206 478 211 490
rect 206 476 207 478
rect 209 476 211 478
rect 206 474 211 476
rect 219 487 223 488
rect 219 485 220 487
rect 222 485 223 487
rect 219 479 223 485
rect 250 487 255 489
rect 219 478 232 479
rect 219 476 224 478
rect 226 476 232 478
rect 219 475 232 476
rect 190 463 191 465
rect 193 464 195 465
rect 193 463 203 464
rect 190 462 203 463
rect 190 460 191 462
rect 193 460 203 462
rect 190 458 203 460
rect 226 470 240 471
rect 226 468 234 470
rect 236 468 240 470
rect 226 467 240 468
rect 250 485 251 487
rect 253 485 255 487
rect 250 483 255 485
rect 250 481 251 483
rect 253 481 255 483
rect 250 480 255 481
rect 250 478 251 480
rect 253 478 255 480
rect 250 476 255 478
rect 226 461 231 467
rect 226 459 228 461
rect 230 459 231 461
rect 226 458 231 459
rect 151 454 175 455
rect 151 452 171 454
rect 173 452 175 454
rect 251 456 255 476
rect 151 451 175 452
rect 243 454 251 456
rect 253 454 255 456
rect 135 450 140 451
rect 243 450 255 454
rect 442 487 458 488
rect 442 485 454 487
rect 456 485 458 487
rect 442 483 458 485
rect 442 455 446 483
rect 490 495 502 496
rect 490 493 498 495
rect 500 493 502 495
rect 490 490 502 493
rect 481 465 486 472
rect 497 478 502 490
rect 497 476 498 478
rect 500 476 502 478
rect 497 474 502 476
rect 510 487 515 489
rect 510 485 512 487
rect 514 485 515 487
rect 510 480 515 485
rect 510 478 512 480
rect 514 478 515 480
rect 510 476 515 478
rect 542 486 546 488
rect 542 484 543 486
rect 545 484 546 486
rect 481 463 482 465
rect 484 464 486 465
rect 484 463 494 464
rect 481 462 494 463
rect 481 460 489 462
rect 491 460 494 462
rect 481 458 494 460
rect 510 462 514 476
rect 510 460 511 462
rect 513 460 514 462
rect 442 454 466 455
rect 442 452 462 454
rect 464 452 466 454
rect 510 456 514 460
rect 542 479 546 484
rect 566 487 570 489
rect 566 485 567 487
rect 569 485 570 487
rect 566 480 570 485
rect 586 487 590 489
rect 586 485 587 487
rect 589 485 590 487
rect 533 478 546 479
rect 533 476 539 478
rect 541 476 546 478
rect 533 475 546 476
rect 554 471 558 480
rect 566 478 567 480
rect 569 479 570 480
rect 586 480 590 485
rect 614 487 630 488
rect 614 486 626 487
rect 614 484 620 486
rect 622 485 626 486
rect 628 485 630 487
rect 622 484 630 485
rect 614 483 630 484
rect 586 479 587 480
rect 569 478 587 479
rect 589 478 590 480
rect 566 476 575 478
rect 577 476 590 478
rect 566 475 590 476
rect 525 470 539 471
rect 525 468 529 470
rect 531 468 536 470
rect 538 468 539 470
rect 525 467 539 468
rect 510 454 512 456
rect 514 454 522 456
rect 442 451 466 452
rect 510 450 522 454
rect 534 458 539 467
rect 554 470 567 471
rect 554 468 558 470
rect 560 468 563 470
rect 565 468 567 470
rect 554 466 567 468
rect 586 461 590 475
rect 594 471 606 472
rect 594 470 603 471
rect 594 468 595 470
rect 597 469 603 470
rect 605 469 606 471
rect 597 468 606 469
rect 594 466 606 468
rect 586 459 587 461
rect 589 459 590 461
rect 586 457 590 459
rect 602 458 606 466
rect 614 455 618 483
rect 662 490 674 496
rect 653 465 658 472
rect 669 478 674 490
rect 669 476 670 478
rect 672 476 674 478
rect 669 474 674 476
rect 653 463 654 465
rect 656 464 658 465
rect 656 463 666 464
rect 653 462 666 463
rect 653 460 663 462
rect 665 460 666 462
rect 653 458 666 460
rect 614 454 638 455
rect 614 452 615 454
rect 617 452 634 454
rect 636 452 638 454
rect 614 451 638 452
rect 27 444 259 445
rect 27 442 33 444
rect 35 442 54 444
rect 56 442 70 444
rect 72 442 82 444
rect 84 442 98 444
rect 100 442 108 444
rect 110 442 153 444
rect 155 442 206 444
rect 208 442 240 444
rect 242 442 250 444
rect 252 442 259 444
rect 27 437 259 442
rect 438 444 678 445
rect 438 442 444 444
rect 446 442 497 444
rect 499 442 513 444
rect 515 442 523 444
rect 525 442 557 444
rect 559 442 616 444
rect 618 442 669 444
rect 671 442 678 444
rect 438 437 678 442
rect 27 432 343 437
rect 27 430 70 432
rect 72 430 80 432
rect 82 430 119 432
rect 121 430 129 432
rect 131 430 190 432
rect 192 430 200 432
rect 202 430 218 432
rect 220 430 230 432
rect 232 430 246 432
rect 248 430 256 432
rect 258 430 290 432
rect 292 430 300 432
rect 302 430 343 432
rect 27 429 343 430
rect 414 432 678 437
rect 414 430 438 432
rect 440 430 448 432
rect 450 430 465 432
rect 467 430 477 432
rect 479 430 511 432
rect 513 430 521 432
rect 523 430 541 432
rect 543 430 551 432
rect 553 430 615 432
rect 617 430 625 432
rect 627 430 678 432
rect 414 429 642 430
rect 644 429 678 430
rect 40 416 44 424
rect 55 422 60 424
rect 55 420 56 422
rect 58 420 60 422
rect 55 418 60 420
rect 28 415 44 416
rect 28 413 29 415
rect 31 413 44 415
rect 28 411 38 413
rect 40 411 44 413
rect 28 410 44 411
rect 56 415 60 418
rect 56 413 57 415
rect 59 413 60 415
rect 48 406 52 408
rect 48 404 49 406
rect 51 404 52 406
rect 48 403 52 404
rect 39 402 52 403
rect 39 400 48 402
rect 50 400 52 402
rect 39 399 52 400
rect 39 395 45 399
rect 56 391 60 413
rect 47 387 60 391
rect 67 420 79 424
rect 67 418 69 420
rect 71 418 79 420
rect 116 420 128 424
rect 67 398 71 418
rect 116 418 118 420
rect 120 418 128 420
rect 91 415 96 416
rect 91 413 92 415
rect 94 413 96 415
rect 91 407 96 413
rect 67 396 72 398
rect 67 394 69 396
rect 71 394 72 396
rect 67 389 72 394
rect 67 387 69 389
rect 71 387 72 389
rect 82 406 96 407
rect 82 404 86 406
rect 88 404 96 406
rect 82 403 96 404
rect 90 398 103 399
rect 90 396 91 398
rect 93 396 96 398
rect 98 396 103 398
rect 90 395 103 396
rect 67 384 72 387
rect 67 382 68 384
rect 70 382 72 384
rect 67 381 72 382
rect 99 386 103 395
rect 116 398 120 418
rect 140 412 145 416
rect 140 410 141 412
rect 143 410 145 412
rect 140 407 145 410
rect 116 396 121 398
rect 116 394 118 396
rect 120 394 121 396
rect 116 393 121 394
rect 116 391 117 393
rect 119 391 121 393
rect 116 389 121 391
rect 116 387 118 389
rect 120 387 121 389
rect 131 406 145 407
rect 131 404 135 406
rect 137 404 145 406
rect 131 403 145 404
rect 176 407 181 416
rect 193 420 205 424
rect 193 418 201 420
rect 203 418 205 420
rect 176 406 190 407
rect 176 404 180 406
rect 182 404 184 406
rect 186 404 190 406
rect 176 403 190 404
rect 139 398 152 399
rect 139 396 145 398
rect 147 396 152 398
rect 139 395 152 396
rect 116 385 121 387
rect 148 389 152 395
rect 148 387 149 389
rect 151 387 152 389
rect 148 386 152 387
rect 169 398 182 399
rect 169 396 174 398
rect 176 396 182 398
rect 169 395 182 396
rect 169 390 173 395
rect 201 401 205 418
rect 201 399 202 401
rect 204 399 205 401
rect 201 398 205 399
rect 169 388 170 390
rect 172 388 173 390
rect 169 386 173 388
rect 200 396 205 398
rect 200 394 201 396
rect 203 394 205 396
rect 200 389 205 394
rect 200 387 201 389
rect 203 387 205 389
rect 200 385 205 387
rect 215 415 219 424
rect 215 413 217 415
rect 215 412 219 413
rect 215 410 216 412
rect 218 410 219 412
rect 215 397 219 410
rect 223 408 227 416
rect 243 420 255 424
rect 243 418 245 420
rect 247 418 255 420
rect 223 406 235 408
rect 223 404 224 406
rect 226 405 235 406
rect 226 404 232 405
rect 223 403 232 404
rect 234 403 235 405
rect 223 402 235 403
rect 215 395 217 397
rect 215 392 219 395
rect 243 398 247 418
rect 287 416 291 424
rect 267 415 272 416
rect 267 413 268 415
rect 270 413 272 415
rect 267 407 272 413
rect 243 396 248 398
rect 243 394 245 396
rect 247 394 248 396
rect 243 393 248 394
rect 215 390 227 392
rect 215 388 217 390
rect 219 388 227 390
rect 215 386 227 388
rect 243 391 244 393
rect 246 391 248 393
rect 243 389 248 391
rect 243 387 245 389
rect 247 387 248 389
rect 258 406 272 407
rect 258 404 262 406
rect 264 404 272 406
rect 258 403 272 404
rect 287 414 289 416
rect 266 398 279 399
rect 266 396 272 398
rect 274 396 276 398
rect 278 396 279 398
rect 266 395 279 396
rect 243 385 248 387
rect 275 386 279 395
rect 287 395 291 414
rect 311 407 315 416
rect 319 415 332 416
rect 319 413 329 415
rect 331 413 332 415
rect 319 410 332 413
rect 302 406 315 407
rect 302 404 306 406
rect 308 404 312 406
rect 314 404 315 406
rect 302 403 315 404
rect 326 406 332 410
rect 326 404 328 406
rect 330 404 332 406
rect 326 403 332 404
rect 424 407 429 416
rect 441 420 453 424
rect 441 418 449 420
rect 451 418 453 420
rect 449 415 453 418
rect 424 406 438 407
rect 424 404 432 406
rect 434 404 435 406
rect 437 404 438 406
rect 424 403 438 404
rect 287 393 289 395
rect 287 391 291 393
rect 310 397 316 399
rect 318 397 332 399
rect 310 395 332 397
rect 417 398 430 399
rect 417 396 422 398
rect 424 396 430 398
rect 417 395 430 396
rect 287 388 300 391
rect 287 386 289 388
rect 291 387 300 388
rect 291 386 292 387
rect 287 382 292 386
rect 287 380 289 382
rect 291 380 292 382
rect 287 378 292 380
rect 318 390 324 395
rect 318 388 321 390
rect 323 388 324 390
rect 318 387 324 388
rect 417 389 421 395
rect 449 413 450 415
rect 452 413 453 415
rect 449 398 453 413
rect 417 387 418 389
rect 420 387 421 389
rect 417 386 421 387
rect 448 396 453 398
rect 448 394 449 396
rect 451 394 453 396
rect 448 389 453 394
rect 448 387 449 389
rect 451 387 453 389
rect 448 385 453 387
rect 462 415 466 424
rect 462 413 464 415
rect 462 397 466 413
rect 470 415 474 416
rect 470 413 471 415
rect 473 413 474 415
rect 497 415 502 416
rect 470 408 474 413
rect 497 413 498 415
rect 500 413 502 415
rect 470 406 482 408
rect 470 404 471 406
rect 473 404 482 406
rect 470 402 482 404
rect 497 407 502 413
rect 514 420 526 424
rect 514 418 522 420
rect 524 418 526 420
rect 497 406 511 407
rect 497 404 505 406
rect 507 404 511 406
rect 497 403 511 404
rect 462 395 464 397
rect 462 392 466 395
rect 490 398 503 399
rect 490 397 495 398
rect 490 395 491 397
rect 493 396 495 397
rect 497 396 503 398
rect 493 395 503 396
rect 462 390 474 392
rect 462 388 464 390
rect 466 389 474 390
rect 466 388 471 389
rect 462 387 471 388
rect 473 387 474 389
rect 462 386 474 387
rect 490 386 494 395
rect 522 398 526 418
rect 521 396 526 398
rect 521 394 522 396
rect 524 394 526 396
rect 521 392 526 394
rect 521 390 523 392
rect 525 390 526 392
rect 521 389 526 390
rect 521 387 522 389
rect 524 387 526 389
rect 521 385 526 387
rect 538 420 550 424
rect 538 418 540 420
rect 542 418 550 420
rect 538 398 542 418
rect 562 407 567 416
rect 538 396 543 398
rect 538 394 540 396
rect 542 394 543 396
rect 538 392 543 394
rect 538 390 540 392
rect 542 390 543 392
rect 538 389 543 390
rect 538 387 540 389
rect 542 387 543 389
rect 553 406 567 407
rect 553 404 554 406
rect 556 404 557 406
rect 559 404 567 406
rect 553 403 567 404
rect 585 410 598 416
rect 585 408 586 410
rect 588 408 591 410
rect 585 406 591 408
rect 585 404 587 406
rect 589 404 591 406
rect 585 403 591 404
rect 602 407 606 416
rect 626 416 630 424
rect 634 423 642 424
rect 634 421 635 423
rect 637 421 642 423
rect 634 420 642 421
rect 665 423 674 424
rect 665 421 667 423
rect 669 421 674 423
rect 665 420 674 421
rect 628 414 630 416
rect 602 406 615 407
rect 602 404 609 406
rect 611 404 612 406
rect 614 404 615 406
rect 602 403 615 404
rect 561 398 574 399
rect 561 396 567 398
rect 569 396 574 398
rect 561 395 574 396
rect 585 397 599 399
rect 601 397 607 399
rect 585 395 607 397
rect 538 385 543 387
rect 570 389 574 395
rect 570 387 571 389
rect 573 387 574 389
rect 570 386 574 387
rect 593 391 599 395
rect 593 389 595 391
rect 597 389 599 391
rect 593 387 599 389
rect 626 395 630 414
rect 638 407 642 420
rect 653 414 666 416
rect 653 412 655 414
rect 657 412 666 414
rect 653 411 666 412
rect 638 406 651 407
rect 638 404 643 406
rect 645 404 651 406
rect 638 403 651 404
rect 662 406 666 411
rect 662 404 663 406
rect 665 404 666 406
rect 662 402 666 404
rect 628 393 630 395
rect 626 391 630 393
rect 617 388 630 391
rect 617 387 626 388
rect 625 386 626 387
rect 628 386 630 388
rect 638 398 657 399
rect 638 396 653 398
rect 655 396 657 398
rect 638 395 657 396
rect 638 389 642 395
rect 670 391 674 420
rect 638 387 639 389
rect 641 387 642 389
rect 638 386 642 387
rect 649 389 674 391
rect 649 387 650 389
rect 652 387 670 389
rect 672 387 674 389
rect 649 386 653 387
rect 625 378 630 386
rect 649 384 650 386
rect 652 384 653 386
rect 649 382 653 384
rect 649 380 650 382
rect 652 380 653 382
rect 649 378 653 380
rect 669 382 674 387
rect 669 380 670 382
rect 672 380 674 382
rect 669 378 674 380
rect 27 372 343 373
rect 27 370 35 372
rect 37 370 43 372
rect 45 370 70 372
rect 72 370 119 372
rect 121 370 200 372
rect 202 370 218 372
rect 220 370 230 372
rect 232 370 246 372
rect 248 370 320 372
rect 322 370 334 372
rect 336 370 343 372
rect 27 365 343 370
rect 414 372 678 373
rect 414 370 448 372
rect 450 370 465 372
rect 467 370 477 372
rect 479 370 521 372
rect 523 370 541 372
rect 543 370 581 372
rect 583 370 595 372
rect 597 370 678 372
rect 414 365 678 370
rect 27 360 291 365
rect 27 358 108 360
rect 110 358 122 360
rect 124 358 162 360
rect 164 358 182 360
rect 184 358 226 360
rect 228 358 238 360
rect 240 358 255 360
rect 257 358 291 360
rect 27 357 291 358
rect 362 360 678 365
rect 362 358 369 360
rect 371 358 383 360
rect 385 358 457 360
rect 459 358 473 360
rect 475 358 485 360
rect 487 358 503 360
rect 505 358 584 360
rect 586 358 633 360
rect 635 358 660 360
rect 662 358 668 360
rect 670 358 678 360
rect 362 357 678 358
rect 31 350 36 352
rect 31 348 33 350
rect 35 348 36 350
rect 31 343 36 348
rect 52 350 56 352
rect 52 348 53 350
rect 55 348 56 350
rect 52 346 56 348
rect 52 344 53 346
rect 55 344 56 346
rect 75 344 80 352
rect 52 343 56 344
rect 31 341 33 343
rect 35 341 53 343
rect 55 341 56 343
rect 31 339 56 341
rect 63 343 67 344
rect 63 341 64 343
rect 66 341 67 343
rect 31 310 35 339
rect 63 335 67 341
rect 48 334 67 335
rect 48 332 50 334
rect 52 332 67 334
rect 48 331 67 332
rect 75 342 77 344
rect 79 343 80 344
rect 79 342 88 343
rect 75 339 88 342
rect 75 337 79 339
rect 75 335 77 337
rect 39 326 43 328
rect 39 324 40 326
rect 42 324 43 326
rect 39 319 43 324
rect 54 326 67 327
rect 54 324 60 326
rect 62 324 67 326
rect 54 323 67 324
rect 39 318 52 319
rect 39 316 48 318
rect 50 316 52 318
rect 39 314 52 316
rect 63 310 67 323
rect 75 316 79 335
rect 106 341 112 343
rect 106 339 108 341
rect 110 339 112 341
rect 106 335 112 339
rect 131 343 135 344
rect 131 341 132 343
rect 134 341 135 343
rect 131 335 135 341
rect 162 343 167 345
rect 98 333 120 335
rect 98 331 104 333
rect 106 331 120 333
rect 131 334 144 335
rect 131 332 136 334
rect 138 332 144 334
rect 131 331 144 332
rect 90 326 103 327
rect 90 324 91 326
rect 93 324 94 326
rect 96 324 103 326
rect 90 323 103 324
rect 75 314 77 316
rect 31 309 40 310
rect 31 307 36 309
rect 38 307 40 309
rect 31 306 40 307
rect 63 309 71 310
rect 63 307 68 309
rect 70 307 71 309
rect 63 306 71 307
rect 75 309 79 314
rect 99 314 103 323
rect 114 326 120 327
rect 114 324 116 326
rect 118 324 120 326
rect 114 322 120 324
rect 114 320 117 322
rect 119 320 120 322
rect 107 314 120 320
rect 138 326 152 327
rect 138 324 146 326
rect 148 324 149 326
rect 151 324 152 326
rect 138 323 152 324
rect 162 341 163 343
rect 165 341 167 343
rect 162 340 167 341
rect 162 338 163 340
rect 165 338 167 340
rect 162 336 167 338
rect 162 334 163 336
rect 165 334 167 336
rect 162 332 167 334
rect 138 314 143 323
rect 75 307 76 309
rect 78 307 79 309
rect 75 306 79 307
rect 163 312 167 332
rect 155 310 163 312
rect 165 310 167 312
rect 155 306 167 310
rect 179 343 184 345
rect 179 341 181 343
rect 183 341 184 343
rect 179 340 184 341
rect 179 338 180 340
rect 182 338 184 340
rect 179 336 184 338
rect 179 334 181 336
rect 183 334 184 336
rect 179 332 184 334
rect 179 312 183 332
rect 211 335 215 344
rect 231 343 243 344
rect 231 341 232 343
rect 234 342 243 343
rect 234 341 239 342
rect 231 340 239 341
rect 241 340 243 342
rect 231 338 243 340
rect 202 334 212 335
rect 202 332 208 334
rect 210 333 212 334
rect 214 333 215 335
rect 210 332 215 333
rect 202 331 215 332
rect 239 335 243 338
rect 241 333 243 335
rect 194 326 208 327
rect 194 324 198 326
rect 200 324 208 326
rect 194 323 208 324
rect 179 310 181 312
rect 183 310 191 312
rect 179 306 191 310
rect 203 317 208 323
rect 223 326 235 328
rect 223 324 232 326
rect 234 324 235 326
rect 223 322 235 324
rect 203 315 205 317
rect 207 315 208 317
rect 231 317 235 322
rect 203 314 208 315
rect 231 315 232 317
rect 234 315 235 317
rect 231 314 235 315
rect 239 317 243 333
rect 241 315 243 317
rect 239 306 243 315
rect 252 343 257 345
rect 252 341 254 343
rect 256 341 257 343
rect 252 336 257 341
rect 252 334 254 336
rect 256 334 257 336
rect 252 332 257 334
rect 284 343 288 344
rect 284 341 285 343
rect 287 341 288 343
rect 252 317 256 332
rect 252 315 253 317
rect 255 315 256 317
rect 284 335 288 341
rect 381 342 387 343
rect 381 340 382 342
rect 384 340 387 342
rect 381 335 387 340
rect 413 350 418 352
rect 413 348 414 350
rect 416 348 418 350
rect 413 344 418 348
rect 413 343 414 344
rect 405 342 414 343
rect 416 342 418 344
rect 405 339 418 342
rect 275 334 288 335
rect 275 332 281 334
rect 283 332 288 334
rect 275 331 288 332
rect 373 333 395 335
rect 373 331 387 333
rect 389 331 395 333
rect 414 337 418 339
rect 416 335 418 337
rect 267 326 281 327
rect 267 324 268 326
rect 270 324 271 326
rect 273 324 281 326
rect 267 323 281 324
rect 252 312 256 315
rect 252 310 254 312
rect 256 310 264 312
rect 252 306 264 310
rect 276 314 281 323
rect 373 326 379 327
rect 373 324 375 326
rect 377 324 379 326
rect 373 320 379 324
rect 390 326 403 327
rect 390 324 391 326
rect 393 324 397 326
rect 399 324 403 326
rect 390 323 403 324
rect 373 317 386 320
rect 373 315 374 317
rect 376 315 386 317
rect 373 314 386 315
rect 390 314 394 323
rect 414 316 418 335
rect 426 335 430 344
rect 457 343 462 345
rect 426 334 439 335
rect 426 332 427 334
rect 429 332 431 334
rect 433 332 439 334
rect 426 331 439 332
rect 416 314 418 316
rect 433 326 447 327
rect 433 324 441 326
rect 443 324 447 326
rect 433 323 447 324
rect 457 341 458 343
rect 460 341 462 343
rect 457 339 462 341
rect 457 337 459 339
rect 461 337 462 339
rect 478 342 490 344
rect 478 340 486 342
rect 488 340 490 342
rect 478 338 490 340
rect 457 336 462 337
rect 457 334 458 336
rect 460 334 462 336
rect 457 332 462 334
rect 433 317 438 323
rect 433 315 435 317
rect 437 315 438 317
rect 433 314 438 315
rect 414 306 418 314
rect 458 312 462 332
rect 486 335 490 338
rect 488 333 490 335
rect 470 327 482 328
rect 470 325 471 327
rect 473 326 482 327
rect 473 325 479 326
rect 470 324 479 325
rect 481 324 482 326
rect 470 322 482 324
rect 450 310 458 312
rect 460 310 462 312
rect 450 306 462 310
rect 478 314 482 322
rect 486 320 490 333
rect 486 318 487 320
rect 489 318 490 320
rect 486 317 490 318
rect 488 315 490 317
rect 486 306 490 315
rect 500 343 505 345
rect 500 341 502 343
rect 504 341 505 343
rect 500 336 505 341
rect 500 334 502 336
rect 504 334 505 336
rect 500 332 505 334
rect 532 342 536 344
rect 532 340 533 342
rect 535 340 536 342
rect 500 331 504 332
rect 500 329 501 331
rect 503 329 504 331
rect 500 312 504 329
rect 532 335 536 340
rect 523 334 536 335
rect 523 332 529 334
rect 531 332 536 334
rect 523 331 536 332
rect 553 343 557 344
rect 553 341 554 343
rect 556 341 557 343
rect 553 335 557 341
rect 584 343 589 345
rect 553 334 566 335
rect 553 332 558 334
rect 560 332 566 334
rect 553 331 566 332
rect 515 326 529 327
rect 515 324 519 326
rect 521 324 523 326
rect 525 324 529 326
rect 515 323 529 324
rect 500 310 502 312
rect 504 310 512 312
rect 500 306 512 310
rect 524 314 529 323
rect 560 326 574 327
rect 560 324 568 326
rect 570 324 574 326
rect 560 323 574 324
rect 584 341 585 343
rect 587 341 589 343
rect 584 339 589 341
rect 584 337 586 339
rect 588 337 589 339
rect 584 336 589 337
rect 584 334 585 336
rect 587 334 589 336
rect 584 332 589 334
rect 560 320 565 323
rect 560 318 562 320
rect 564 318 565 320
rect 560 314 565 318
rect 585 312 589 332
rect 602 335 606 344
rect 633 348 638 349
rect 633 346 635 348
rect 637 346 638 348
rect 633 343 638 346
rect 602 334 615 335
rect 602 332 607 334
rect 609 332 612 334
rect 614 332 615 334
rect 602 331 615 332
rect 609 326 623 327
rect 609 324 617 326
rect 619 324 623 326
rect 609 323 623 324
rect 633 341 634 343
rect 636 341 638 343
rect 633 336 638 341
rect 633 334 634 336
rect 636 334 638 336
rect 633 332 638 334
rect 609 317 614 323
rect 609 315 611 317
rect 613 315 614 317
rect 609 314 614 315
rect 577 310 585 312
rect 587 310 589 312
rect 634 312 638 332
rect 577 306 589 310
rect 626 310 634 312
rect 636 310 638 312
rect 626 306 638 310
rect 645 339 658 343
rect 645 317 649 339
rect 660 331 666 335
rect 653 330 666 331
rect 653 328 655 330
rect 657 328 666 330
rect 653 327 666 328
rect 653 326 657 327
rect 653 324 654 326
rect 656 324 657 326
rect 653 322 657 324
rect 645 315 646 317
rect 648 315 649 317
rect 645 312 649 315
rect 661 319 677 320
rect 661 317 665 319
rect 667 317 677 319
rect 661 315 674 317
rect 676 315 677 317
rect 661 314 677 315
rect 645 310 650 312
rect 645 308 647 310
rect 649 308 650 310
rect 645 306 650 308
rect 661 306 665 314
rect 27 300 61 301
rect 63 300 291 301
rect 27 298 78 300
rect 80 298 88 300
rect 90 298 152 300
rect 154 298 162 300
rect 164 298 182 300
rect 184 298 192 300
rect 194 298 226 300
rect 228 298 238 300
rect 240 298 255 300
rect 257 298 265 300
rect 267 298 291 300
rect 27 293 291 298
rect 362 300 678 301
rect 362 298 403 300
rect 405 298 413 300
rect 415 298 447 300
rect 449 298 457 300
rect 459 298 473 300
rect 475 298 485 300
rect 487 298 503 300
rect 505 298 513 300
rect 515 298 574 300
rect 576 298 584 300
rect 586 298 623 300
rect 625 298 633 300
rect 635 298 678 300
rect 362 293 678 298
rect 27 288 295 293
rect 27 286 34 288
rect 36 286 87 288
rect 89 286 146 288
rect 148 286 180 288
rect 182 286 190 288
rect 192 286 206 288
rect 208 286 259 288
rect 261 286 274 288
rect 276 286 286 288
rect 288 286 295 288
rect 27 285 295 286
rect 446 288 678 293
rect 446 286 453 288
rect 455 286 463 288
rect 465 286 497 288
rect 499 286 550 288
rect 552 286 595 288
rect 597 286 605 288
rect 607 286 621 288
rect 623 286 633 288
rect 635 286 649 288
rect 651 286 670 288
rect 672 286 678 288
rect 446 285 678 286
rect 67 278 91 279
rect 67 276 69 278
rect 71 276 88 278
rect 90 276 91 278
rect 67 275 91 276
rect 39 270 52 272
rect 39 268 40 270
rect 42 268 52 270
rect 39 267 52 268
rect 39 266 49 267
rect 47 265 49 266
rect 51 265 52 267
rect 31 254 36 256
rect 31 252 33 254
rect 35 252 36 254
rect 31 240 36 252
rect 47 258 52 265
rect 31 234 43 240
rect 87 247 91 275
rect 99 264 103 272
rect 115 271 119 273
rect 115 269 116 271
rect 118 269 119 271
rect 99 262 111 264
rect 99 261 108 262
rect 99 259 100 261
rect 102 260 108 261
rect 110 260 111 262
rect 102 259 111 260
rect 99 258 111 259
rect 115 255 119 269
rect 138 262 151 264
rect 138 260 140 262
rect 142 260 145 262
rect 147 260 151 262
rect 138 259 151 260
rect 166 263 171 272
rect 183 276 195 280
rect 239 278 263 279
rect 183 274 191 276
rect 193 274 195 276
rect 166 262 180 263
rect 166 260 167 262
rect 169 260 174 262
rect 176 260 180 262
rect 166 259 180 260
rect 115 254 139 255
rect 115 252 128 254
rect 130 252 139 254
rect 115 250 116 252
rect 118 251 136 252
rect 118 250 119 251
rect 75 246 91 247
rect 75 245 83 246
rect 75 243 77 245
rect 79 244 83 245
rect 85 244 91 246
rect 79 243 91 244
rect 75 242 91 243
rect 115 245 119 250
rect 135 250 136 251
rect 138 250 139 252
rect 147 250 151 259
rect 159 254 172 255
rect 159 252 164 254
rect 166 252 172 254
rect 159 251 172 252
rect 115 243 116 245
rect 118 243 119 245
rect 115 241 119 243
rect 135 245 139 250
rect 135 243 136 245
rect 138 243 139 245
rect 135 241 139 243
rect 159 246 163 251
rect 191 270 195 274
rect 239 276 241 278
rect 243 276 263 278
rect 239 275 263 276
rect 191 268 192 270
rect 194 268 195 270
rect 191 254 195 268
rect 211 270 224 272
rect 211 268 214 270
rect 216 268 224 270
rect 211 267 224 268
rect 211 266 221 267
rect 219 265 221 266
rect 223 265 224 267
rect 159 244 160 246
rect 162 244 163 246
rect 159 242 163 244
rect 190 252 195 254
rect 190 250 191 252
rect 193 250 195 252
rect 190 245 195 250
rect 190 243 191 245
rect 193 243 195 245
rect 190 241 195 243
rect 203 254 208 256
rect 203 252 205 254
rect 207 252 208 254
rect 203 240 208 252
rect 219 258 224 265
rect 203 237 215 240
rect 203 235 205 237
rect 207 235 215 237
rect 203 234 215 235
rect 259 247 263 275
rect 247 245 263 247
rect 247 243 249 245
rect 251 243 263 245
rect 247 242 263 243
rect 271 271 275 280
rect 271 269 273 271
rect 271 253 275 269
rect 279 270 283 272
rect 450 276 462 280
rect 565 279 570 280
rect 450 274 452 276
rect 454 274 462 276
rect 530 278 554 279
rect 279 268 280 270
rect 282 268 283 270
rect 279 264 283 268
rect 279 262 291 264
rect 279 260 280 262
rect 282 260 291 262
rect 279 258 291 260
rect 271 251 273 253
rect 271 248 275 251
rect 450 254 454 274
rect 530 276 532 278
rect 534 276 554 278
rect 530 275 554 276
rect 474 271 479 272
rect 474 269 475 271
rect 477 269 479 271
rect 474 263 479 269
rect 450 252 455 254
rect 450 250 452 252
rect 454 250 455 252
rect 450 249 455 250
rect 271 246 283 248
rect 271 244 273 246
rect 275 244 280 246
rect 282 244 283 246
rect 271 242 283 244
rect 450 247 452 249
rect 454 247 455 249
rect 450 245 455 247
rect 450 243 452 245
rect 454 243 455 245
rect 465 262 479 263
rect 465 260 469 262
rect 471 260 479 262
rect 465 259 479 260
rect 502 270 515 272
rect 502 268 512 270
rect 514 268 515 270
rect 502 267 515 268
rect 502 266 512 267
rect 510 265 512 266
rect 514 265 515 267
rect 473 254 486 255
rect 473 252 479 254
rect 481 252 486 254
rect 473 251 486 252
rect 450 241 455 243
rect 482 245 486 251
rect 482 243 483 245
rect 485 243 486 245
rect 482 242 486 243
rect 494 254 499 256
rect 494 252 496 254
rect 498 252 499 254
rect 494 240 499 252
rect 510 258 515 265
rect 494 238 506 240
rect 494 236 503 238
rect 505 236 506 238
rect 494 234 506 236
rect 550 247 554 275
rect 565 277 567 279
rect 569 277 570 279
rect 565 272 570 277
rect 565 267 586 272
rect 598 276 610 280
rect 598 274 606 276
rect 608 274 610 276
rect 581 263 586 267
rect 581 262 595 263
rect 581 260 589 262
rect 591 260 595 262
rect 581 259 595 260
rect 538 245 554 247
rect 538 243 540 245
rect 542 243 554 245
rect 538 242 554 243
rect 574 254 587 255
rect 574 252 579 254
rect 581 252 587 254
rect 574 251 587 252
rect 574 246 578 251
rect 606 270 610 274
rect 634 279 638 280
rect 634 277 635 279
rect 637 277 638 279
rect 626 271 630 272
rect 606 268 607 270
rect 609 268 610 270
rect 606 254 610 268
rect 626 269 627 271
rect 629 269 630 271
rect 626 264 630 269
rect 634 271 638 277
rect 655 279 677 280
rect 655 277 659 279
rect 661 277 674 279
rect 676 277 677 279
rect 655 276 677 277
rect 662 274 674 276
rect 636 269 638 271
rect 618 262 630 264
rect 618 260 627 262
rect 629 260 630 262
rect 618 258 630 260
rect 574 244 575 246
rect 577 244 578 246
rect 574 242 578 244
rect 605 252 610 254
rect 605 250 606 252
rect 608 250 610 252
rect 605 245 610 250
rect 634 253 638 269
rect 654 266 658 272
rect 646 265 658 266
rect 646 263 653 265
rect 655 263 658 265
rect 670 271 674 274
rect 670 269 671 271
rect 673 269 674 271
rect 646 262 658 263
rect 662 262 666 264
rect 646 261 650 262
rect 646 259 647 261
rect 649 259 650 261
rect 646 258 650 259
rect 662 260 663 262
rect 665 260 666 262
rect 662 258 666 260
rect 654 254 666 258
rect 636 251 638 253
rect 634 248 638 251
rect 646 253 658 254
rect 646 251 647 253
rect 649 251 658 253
rect 646 250 658 251
rect 605 243 606 245
rect 608 243 610 245
rect 605 241 610 243
rect 626 246 638 248
rect 670 246 674 269
rect 626 244 634 246
rect 636 244 638 246
rect 626 242 638 244
rect 665 245 674 246
rect 665 243 667 245
rect 669 243 674 245
rect 665 242 674 243
rect 665 238 671 242
rect 665 236 667 238
rect 669 236 671 238
rect 665 235 671 236
rect 27 228 295 229
rect 27 226 67 228
rect 69 226 138 228
rect 140 226 146 228
rect 148 226 190 228
rect 192 226 239 228
rect 241 226 274 228
rect 276 226 286 228
rect 288 226 295 228
rect 27 221 295 226
rect 446 228 678 229
rect 446 226 453 228
rect 455 226 530 228
rect 532 226 605 228
rect 607 226 621 228
rect 623 226 633 228
rect 635 226 678 228
rect 27 216 203 221
rect 27 214 84 216
rect 86 214 96 216
rect 98 214 114 216
rect 116 214 203 216
rect 27 213 203 214
rect 446 216 678 226
rect 446 214 479 216
rect 481 214 493 216
rect 495 214 636 216
rect 638 214 678 216
rect 446 213 678 214
rect 47 199 53 201
rect 47 197 50 199
rect 52 197 53 199
rect 47 195 53 197
rect 47 193 48 195
rect 50 193 53 195
rect 89 198 101 200
rect 111 199 116 201
rect 89 196 97 198
rect 99 196 101 198
rect 89 194 101 196
rect 108 198 113 199
rect 108 196 109 198
rect 111 197 113 198
rect 115 197 116 199
rect 111 196 116 197
rect 108 195 116 196
rect 47 192 53 193
rect 47 191 50 192
rect 31 190 50 191
rect 52 190 53 192
rect 31 187 53 190
rect 63 191 68 192
rect 63 189 65 191
rect 67 189 68 191
rect 31 167 35 187
rect 63 183 68 189
rect 97 192 98 194
rect 100 192 101 194
rect 97 191 101 192
rect 99 189 101 191
rect 51 182 68 183
rect 51 180 53 182
rect 55 180 68 182
rect 51 179 68 180
rect 81 182 93 184
rect 81 180 84 182
rect 86 180 90 182
rect 92 180 93 182
rect 41 177 45 179
rect 81 178 93 180
rect 41 175 42 177
rect 44 175 45 177
rect 41 174 68 175
rect 41 172 57 174
rect 59 172 64 174
rect 66 172 68 174
rect 41 171 68 172
rect 31 166 49 167
rect 31 164 45 166
rect 47 164 49 166
rect 31 163 49 164
rect 63 162 68 171
rect 89 170 93 178
rect 97 173 101 189
rect 99 171 101 173
rect 97 162 101 171
rect 111 192 116 195
rect 111 190 113 192
rect 115 190 116 192
rect 111 188 116 190
rect 111 168 115 188
rect 143 191 147 200
rect 171 199 177 201
rect 171 197 174 199
rect 176 197 177 199
rect 171 196 177 197
rect 171 194 174 196
rect 176 194 177 196
rect 171 192 177 194
rect 446 200 451 208
rect 446 198 448 200
rect 450 199 451 200
rect 450 198 459 199
rect 446 195 459 198
rect 446 193 450 195
rect 171 191 174 192
rect 134 190 147 191
rect 134 188 140 190
rect 142 188 144 190
rect 146 188 147 190
rect 134 187 147 188
rect 155 190 174 191
rect 176 190 177 192
rect 155 187 177 190
rect 126 182 140 183
rect 126 180 130 182
rect 132 180 140 182
rect 126 179 140 180
rect 111 166 113 168
rect 115 166 123 168
rect 111 162 123 166
rect 135 174 140 179
rect 135 172 136 174
rect 138 172 140 174
rect 135 170 140 172
rect 155 167 159 187
rect 187 183 192 192
rect 446 191 448 193
rect 175 182 219 183
rect 175 180 177 182
rect 179 180 216 182
rect 218 180 219 182
rect 175 179 219 180
rect 165 177 169 179
rect 165 175 166 177
rect 168 175 169 177
rect 165 174 192 175
rect 165 172 166 174
rect 168 172 188 174
rect 190 172 192 174
rect 165 171 192 172
rect 155 166 173 167
rect 155 164 169 166
rect 171 164 173 166
rect 155 163 173 164
rect 187 162 192 171
rect 446 172 450 191
rect 477 198 483 199
rect 477 196 480 198
rect 482 196 483 198
rect 477 191 483 196
rect 594 199 606 200
rect 506 198 534 199
rect 506 196 507 198
rect 509 197 534 198
rect 536 197 543 199
rect 509 196 543 197
rect 506 195 543 196
rect 594 197 603 199
rect 605 197 606 199
rect 469 189 491 191
rect 469 187 475 189
rect 477 187 491 189
rect 461 182 474 183
rect 461 180 462 182
rect 464 180 465 182
rect 467 180 474 182
rect 461 179 474 180
rect 446 170 448 172
rect 446 166 450 170
rect 470 170 474 179
rect 485 182 491 183
rect 485 180 487 182
rect 489 180 491 182
rect 485 176 491 180
rect 478 174 491 176
rect 478 172 479 174
rect 481 172 491 174
rect 478 170 491 172
rect 446 164 447 166
rect 449 164 450 166
rect 446 162 450 164
rect 506 166 510 195
rect 594 194 606 197
rect 578 191 590 192
rect 514 190 559 191
rect 514 188 515 190
rect 517 188 559 190
rect 514 187 559 188
rect 514 174 518 187
rect 555 183 559 187
rect 578 189 584 191
rect 586 189 590 191
rect 578 186 590 189
rect 578 184 580 186
rect 514 172 515 174
rect 517 172 518 174
rect 514 170 518 172
rect 522 179 551 183
rect 555 182 562 183
rect 555 180 558 182
rect 560 180 562 182
rect 555 179 562 180
rect 522 174 528 179
rect 547 176 551 179
rect 578 178 582 184
rect 594 182 598 184
rect 594 180 595 182
rect 597 180 598 182
rect 594 176 598 180
rect 522 172 525 174
rect 527 172 528 174
rect 522 170 528 172
rect 535 174 543 175
rect 535 172 537 174
rect 539 172 543 174
rect 535 171 543 172
rect 547 174 548 176
rect 550 175 551 176
rect 586 175 598 176
rect 550 174 559 175
rect 547 172 556 174
rect 558 172 559 174
rect 547 171 559 172
rect 586 173 591 175
rect 593 173 598 175
rect 538 167 543 171
rect 586 170 598 173
rect 538 166 551 167
rect 506 165 534 166
rect 506 163 508 165
rect 510 163 530 165
rect 532 163 534 165
rect 506 162 534 163
rect 538 164 548 166
rect 550 164 551 166
rect 538 162 551 164
rect 602 166 606 194
rect 597 165 606 166
rect 597 163 599 165
rect 601 163 606 165
rect 614 199 630 200
rect 614 197 626 199
rect 628 197 630 199
rect 614 195 630 197
rect 614 175 618 195
rect 662 202 674 208
rect 614 173 615 175
rect 617 173 618 175
rect 614 167 618 173
rect 653 177 658 184
rect 669 190 674 202
rect 669 188 670 190
rect 672 188 674 190
rect 669 186 674 188
rect 653 175 654 177
rect 656 176 658 177
rect 656 175 666 176
rect 653 174 666 175
rect 653 172 663 174
rect 665 172 666 174
rect 653 170 666 172
rect 614 166 638 167
rect 614 164 634 166
rect 636 164 638 166
rect 614 163 638 164
rect 597 162 606 163
rect 27 156 203 157
rect 27 154 70 156
rect 72 154 84 156
rect 86 154 96 156
rect 98 154 114 156
rect 116 154 124 156
rect 126 154 194 156
rect 196 154 203 156
rect 27 149 203 154
rect 446 156 678 157
rect 446 154 449 156
rect 451 154 459 156
rect 461 154 519 156
rect 521 154 541 156
rect 543 154 557 156
rect 559 154 616 156
rect 618 154 669 156
rect 671 154 678 156
rect 446 149 678 154
rect 27 144 211 149
rect 27 142 34 144
rect 36 142 87 144
rect 89 142 158 144
rect 160 142 168 144
rect 170 142 188 144
rect 190 142 200 144
rect 202 142 211 144
rect 27 141 211 142
rect 418 144 678 149
rect 418 142 429 144
rect 431 142 473 144
rect 475 142 551 144
rect 553 142 561 144
rect 563 142 595 144
rect 597 142 605 144
rect 607 142 621 144
rect 623 142 633 144
rect 635 142 678 144
rect 418 141 678 142
rect 99 135 108 136
rect 67 134 91 135
rect 67 132 69 134
rect 71 132 91 134
rect 67 131 91 132
rect 39 127 52 128
rect 39 125 40 127
rect 42 125 52 127
rect 39 123 52 125
rect 39 122 49 123
rect 47 121 49 122
rect 51 121 52 123
rect 31 110 36 112
rect 31 108 33 110
rect 35 108 36 110
rect 31 96 36 108
rect 47 114 52 121
rect 87 126 91 131
rect 87 124 88 126
rect 90 124 91 126
rect 31 90 43 96
rect 87 103 91 124
rect 75 101 91 103
rect 75 99 77 101
rect 79 99 81 101
rect 83 99 91 101
rect 75 98 91 99
rect 99 133 100 135
rect 102 133 104 135
rect 106 133 108 135
rect 99 132 108 133
rect 99 104 103 132
rect 107 126 119 128
rect 107 124 108 126
rect 110 124 119 126
rect 107 122 119 124
rect 144 127 149 128
rect 144 125 145 127
rect 147 125 149 127
rect 107 118 111 122
rect 107 116 108 118
rect 110 116 111 118
rect 107 114 111 116
rect 123 114 127 120
rect 144 119 149 125
rect 161 132 173 136
rect 161 130 169 132
rect 171 130 173 132
rect 144 118 158 119
rect 144 116 152 118
rect 154 116 158 118
rect 144 115 158 116
rect 125 112 127 114
rect 115 109 127 112
rect 115 107 117 109
rect 119 107 127 109
rect 115 106 127 107
rect 137 110 150 111
rect 137 108 142 110
rect 144 108 150 110
rect 137 107 150 108
rect 99 98 111 104
rect 137 101 141 107
rect 169 112 173 130
rect 169 110 170 112
rect 172 110 173 112
rect 137 99 138 101
rect 140 99 141 101
rect 137 98 141 99
rect 168 108 173 110
rect 168 106 169 108
rect 171 106 173 108
rect 168 101 173 106
rect 168 99 169 101
rect 171 99 173 101
rect 168 97 173 99
rect 185 127 189 136
rect 185 125 187 127
rect 185 109 189 125
rect 193 120 197 128
rect 430 134 442 136
rect 430 132 439 134
rect 441 132 442 134
rect 430 130 442 132
rect 460 135 490 136
rect 460 133 462 135
rect 464 133 484 135
rect 486 133 490 135
rect 460 131 490 133
rect 430 125 434 130
rect 447 126 472 127
rect 430 123 431 125
rect 433 123 434 125
rect 430 122 434 123
rect 438 123 442 125
rect 447 124 449 126
rect 451 124 454 126
rect 456 124 468 126
rect 470 124 472 126
rect 447 123 472 124
rect 478 124 482 126
rect 438 121 439 123
rect 441 121 442 123
rect 193 119 205 120
rect 193 118 198 119
rect 193 116 194 118
rect 196 117 198 118
rect 200 117 205 119
rect 438 119 442 121
rect 196 116 205 117
rect 193 114 205 116
rect 427 117 433 118
rect 427 115 429 117
rect 431 115 433 117
rect 438 115 451 119
rect 461 115 467 123
rect 478 122 479 124
rect 481 122 482 124
rect 427 111 433 115
rect 447 111 451 115
rect 478 111 482 122
rect 185 107 187 109
rect 185 104 189 107
rect 427 107 442 111
rect 447 110 482 111
rect 447 108 479 110
rect 481 108 482 110
rect 447 107 482 108
rect 185 102 197 104
rect 185 100 187 102
rect 189 100 190 102
rect 192 100 197 102
rect 185 98 197 100
rect 438 95 442 107
rect 486 103 490 131
rect 521 127 534 128
rect 521 125 522 127
rect 524 125 534 127
rect 521 122 534 125
rect 538 127 542 128
rect 538 125 539 127
rect 541 125 542 127
rect 494 117 498 119
rect 496 115 498 117
rect 521 118 527 122
rect 521 116 523 118
rect 525 116 527 118
rect 521 115 527 116
rect 538 119 542 125
rect 562 128 566 136
rect 564 126 566 128
rect 538 118 551 119
rect 538 116 545 118
rect 547 116 551 118
rect 538 115 551 116
rect 457 102 490 103
rect 457 100 459 102
rect 461 100 487 102
rect 489 100 490 102
rect 457 99 490 100
rect 494 95 498 115
rect 521 110 535 111
rect 521 108 531 110
rect 533 109 535 110
rect 537 109 543 111
rect 533 108 543 109
rect 521 107 543 108
rect 438 94 498 95
rect 438 92 495 94
rect 497 92 498 94
rect 438 91 498 92
rect 529 99 535 107
rect 562 107 566 126
rect 581 124 586 128
rect 581 122 583 124
rect 585 122 586 124
rect 598 132 610 136
rect 598 130 606 132
rect 608 130 610 132
rect 581 119 586 122
rect 581 118 595 119
rect 581 116 589 118
rect 591 116 595 118
rect 581 115 595 116
rect 564 105 566 107
rect 562 103 566 105
rect 553 102 566 103
rect 553 100 554 102
rect 556 100 566 102
rect 553 99 562 100
rect 561 98 562 99
rect 564 98 566 100
rect 574 110 587 111
rect 574 108 579 110
rect 581 108 584 110
rect 586 108 587 110
rect 574 107 587 108
rect 574 98 578 107
rect 606 110 610 130
rect 634 135 638 136
rect 634 133 635 135
rect 637 133 638 135
rect 626 120 630 128
rect 634 127 638 133
rect 665 135 674 136
rect 665 133 667 135
rect 669 133 674 135
rect 665 132 674 133
rect 636 125 638 127
rect 618 118 630 120
rect 618 117 627 118
rect 618 115 619 117
rect 621 116 627 117
rect 629 116 630 118
rect 621 115 630 116
rect 618 114 630 115
rect 605 108 610 110
rect 605 106 606 108
rect 608 106 610 108
rect 605 104 610 106
rect 634 109 638 125
rect 654 127 666 128
rect 654 125 655 127
rect 657 125 666 127
rect 654 122 666 125
rect 636 107 638 109
rect 634 104 638 107
rect 646 114 650 120
rect 662 118 666 122
rect 662 116 663 118
rect 665 116 666 118
rect 646 112 648 114
rect 662 114 666 116
rect 670 125 674 132
rect 670 123 671 125
rect 673 123 674 125
rect 646 109 658 112
rect 646 107 647 109
rect 649 107 658 109
rect 646 106 658 107
rect 670 104 674 123
rect 605 102 607 104
rect 609 102 610 104
rect 605 101 610 102
rect 561 90 566 98
rect 605 99 606 101
rect 608 99 610 101
rect 605 97 610 99
rect 626 102 638 104
rect 626 100 634 102
rect 636 100 638 102
rect 626 98 638 100
rect 662 98 674 104
rect 27 84 211 85
rect 27 82 67 84
rect 69 82 168 84
rect 170 82 188 84
rect 190 82 200 84
rect 202 82 211 84
rect 27 72 211 82
rect 418 84 678 85
rect 418 82 429 84
rect 431 82 451 84
rect 453 82 491 84
rect 493 82 517 84
rect 519 82 531 84
rect 533 82 605 84
rect 607 82 621 84
rect 623 82 633 84
rect 635 82 678 84
rect 418 77 678 82
rect 27 70 82 72
rect 84 70 94 72
rect 96 70 132 72
rect 134 70 184 72
rect 186 70 211 72
rect 27 69 211 70
rect 369 72 678 77
rect 369 70 379 72
rect 381 70 391 72
rect 393 70 411 72
rect 413 70 488 72
rect 490 70 565 72
rect 567 70 636 72
rect 638 70 678 72
rect 369 69 678 70
rect 47 55 53 57
rect 47 53 50 55
rect 52 53 53 55
rect 47 48 53 53
rect 87 54 99 56
rect 87 53 95 54
rect 87 51 90 53
rect 92 52 95 53
rect 97 52 99 54
rect 92 51 99 52
rect 87 50 99 51
rect 47 47 50 48
rect 31 46 50 47
rect 52 46 53 48
rect 31 44 32 46
rect 34 44 53 46
rect 31 43 53 44
rect 63 47 68 48
rect 63 45 65 47
rect 67 45 68 47
rect 31 23 35 43
rect 63 39 68 45
rect 95 47 99 50
rect 97 45 99 47
rect 51 38 68 39
rect 51 36 53 38
rect 55 36 68 38
rect 51 35 68 36
rect 79 38 91 40
rect 79 36 88 38
rect 90 36 91 38
rect 41 33 45 35
rect 79 34 91 36
rect 41 31 42 33
rect 44 31 45 33
rect 41 30 68 31
rect 41 28 42 30
rect 44 28 64 30
rect 66 28 68 30
rect 87 29 91 34
rect 41 27 68 28
rect 31 22 49 23
rect 31 20 42 22
rect 44 20 45 22
rect 47 20 49 22
rect 31 19 49 20
rect 63 18 68 27
rect 87 27 88 29
rect 90 27 91 29
rect 87 26 91 27
rect 95 29 99 45
rect 97 27 99 29
rect 95 18 99 27
rect 110 55 126 56
rect 110 53 122 55
rect 124 53 126 55
rect 110 51 126 53
rect 110 23 114 51
rect 158 63 170 64
rect 158 61 167 63
rect 169 61 170 63
rect 158 58 170 61
rect 149 39 154 40
rect 149 37 151 39
rect 153 37 154 39
rect 149 33 154 37
rect 165 46 170 58
rect 384 55 396 56
rect 191 54 208 55
rect 191 52 193 54
rect 195 52 198 54
rect 200 52 208 54
rect 191 51 208 52
rect 165 44 166 46
rect 168 44 170 46
rect 165 42 170 44
rect 180 46 193 47
rect 180 44 190 46
rect 192 44 193 46
rect 180 43 193 44
rect 180 39 184 43
rect 149 31 150 33
rect 152 32 154 33
rect 152 31 162 32
rect 149 26 162 31
rect 180 37 182 39
rect 180 34 184 37
rect 204 32 208 51
rect 384 53 385 55
rect 387 54 396 55
rect 387 53 392 54
rect 384 52 392 53
rect 394 52 396 54
rect 384 50 396 52
rect 392 47 396 50
rect 394 45 396 47
rect 376 38 388 40
rect 376 37 385 38
rect 376 35 378 37
rect 380 36 385 37
rect 387 36 388 38
rect 380 35 388 36
rect 376 34 388 35
rect 188 29 208 32
rect 188 27 193 29
rect 195 27 208 29
rect 188 26 208 27
rect 384 26 388 34
rect 110 22 134 23
rect 110 20 130 22
rect 132 20 134 22
rect 392 29 396 45
rect 412 48 416 64
rect 420 62 425 64
rect 420 60 422 62
rect 424 60 425 62
rect 420 56 425 60
rect 420 55 456 56
rect 420 53 422 55
rect 424 53 442 55
rect 444 53 456 55
rect 420 52 456 53
rect 444 50 456 52
rect 412 47 424 48
rect 412 45 413 47
rect 415 45 424 47
rect 412 44 424 45
rect 394 27 396 29
rect 110 19 134 20
rect 392 18 396 27
rect 412 38 416 40
rect 412 36 413 38
rect 415 36 416 38
rect 412 32 416 36
rect 420 34 424 44
rect 434 45 440 48
rect 434 43 435 45
rect 437 43 440 45
rect 434 38 440 43
rect 428 34 440 38
rect 444 38 448 40
rect 444 36 445 38
rect 447 36 448 38
rect 444 35 448 36
rect 412 30 413 32
rect 415 30 416 32
rect 412 24 416 30
rect 428 29 432 34
rect 444 33 445 35
rect 447 33 448 35
rect 444 30 448 33
rect 428 27 429 29
rect 431 27 432 29
rect 412 18 424 24
rect 428 18 432 27
rect 436 26 448 30
rect 436 18 440 26
rect 452 22 456 50
rect 444 21 456 22
rect 444 19 446 21
rect 448 19 453 21
rect 455 19 456 21
rect 466 55 482 56
rect 466 53 478 55
rect 480 53 482 55
rect 466 51 482 53
rect 466 23 470 51
rect 514 63 526 64
rect 514 61 517 63
rect 519 61 526 63
rect 514 58 526 61
rect 505 33 510 40
rect 521 46 526 58
rect 521 44 522 46
rect 524 44 526 46
rect 521 42 526 44
rect 534 55 538 56
rect 534 53 535 55
rect 537 53 538 55
rect 534 47 538 53
rect 597 62 603 63
rect 597 60 599 62
rect 601 60 603 62
rect 597 59 603 60
rect 597 57 598 59
rect 600 57 603 59
rect 565 55 570 57
rect 534 46 547 47
rect 534 44 539 46
rect 541 44 547 46
rect 534 43 547 44
rect 505 31 506 33
rect 508 32 510 33
rect 508 31 518 32
rect 505 29 518 31
rect 505 27 515 29
rect 517 27 518 29
rect 505 26 518 27
rect 541 38 555 39
rect 541 36 549 38
rect 551 36 555 38
rect 541 35 555 36
rect 565 53 566 55
rect 568 53 570 55
rect 565 48 570 53
rect 597 56 603 57
rect 597 55 606 56
rect 597 53 599 55
rect 601 53 606 55
rect 597 52 606 53
rect 565 46 566 48
rect 568 46 570 48
rect 565 44 570 46
rect 541 32 546 35
rect 541 30 542 32
rect 544 30 546 32
rect 541 26 546 30
rect 466 22 490 23
rect 466 20 486 22
rect 488 20 490 22
rect 566 24 570 44
rect 586 46 590 48
rect 586 44 587 46
rect 589 44 590 46
rect 586 40 598 44
rect 578 36 582 40
rect 594 38 598 40
rect 594 36 595 38
rect 597 36 598 38
rect 578 35 590 36
rect 578 33 585 35
rect 587 33 590 35
rect 594 34 598 36
rect 578 32 590 33
rect 586 29 590 32
rect 586 27 587 29
rect 589 27 590 29
rect 586 26 590 27
rect 466 19 490 20
rect 558 23 566 24
rect 558 21 559 23
rect 561 22 566 23
rect 568 22 570 24
rect 561 21 570 22
rect 444 18 456 19
rect 558 18 570 21
rect 602 24 606 52
rect 594 22 606 24
rect 589 21 606 22
rect 589 19 591 21
rect 593 19 606 21
rect 614 55 630 56
rect 614 54 626 55
rect 614 52 619 54
rect 621 53 626 54
rect 628 53 630 55
rect 621 52 630 53
rect 614 51 630 52
rect 614 29 618 51
rect 662 58 674 64
rect 614 27 615 29
rect 617 27 618 29
rect 653 33 658 40
rect 669 46 674 58
rect 669 44 670 46
rect 672 44 674 46
rect 669 42 674 44
rect 653 31 654 33
rect 656 32 658 33
rect 656 31 666 32
rect 614 23 618 27
rect 653 30 666 31
rect 653 28 663 30
rect 665 28 666 30
rect 653 26 666 28
rect 614 22 638 23
rect 614 20 634 22
rect 636 20 638 22
rect 614 19 638 20
rect 589 18 606 19
rect 27 12 211 13
rect 27 10 70 12
rect 72 10 82 12
rect 84 10 94 12
rect 96 10 112 12
rect 114 10 165 12
rect 167 10 183 12
rect 185 10 203 12
rect 205 10 211 12
rect 27 5 211 10
rect 369 12 678 13
rect 369 10 379 12
rect 381 10 391 12
rect 393 10 414 12
rect 416 10 468 12
rect 470 10 521 12
rect 523 10 555 12
rect 557 10 565 12
rect 567 10 581 12
rect 583 10 602 12
rect 604 10 616 12
rect 618 10 669 12
rect 671 10 678 12
rect 369 5 678 10
<< alu2 >>
rect 249 711 328 712
rect 143 709 191 710
rect 143 707 144 709
rect 146 707 191 709
rect 249 709 250 711
rect 252 709 328 711
rect 249 708 328 709
rect 143 706 191 707
rect 39 702 43 704
rect 39 700 40 702
rect 42 700 43 702
rect 87 703 119 704
rect 87 701 88 703
rect 90 701 116 703
rect 118 701 119 703
rect 187 703 191 706
rect 187 701 188 703
rect 190 701 191 703
rect 87 700 119 701
rect 160 700 164 701
rect 187 700 191 701
rect 265 703 277 704
rect 265 701 266 703
rect 268 701 274 703
rect 276 701 277 703
rect 265 700 277 701
rect 289 700 302 701
rect 31 607 35 608
rect 31 605 32 607
rect 34 605 35 607
rect 31 592 35 605
rect 31 590 32 592
rect 34 590 35 592
rect 31 589 35 590
rect 39 558 43 700
rect 160 698 161 700
rect 163 698 164 700
rect 289 698 290 700
rect 292 698 299 700
rect 301 698 302 700
rect 160 696 164 698
rect 160 694 161 696
rect 163 694 164 696
rect 160 693 164 694
rect 257 697 261 698
rect 289 697 302 698
rect 257 695 258 697
rect 260 695 261 697
rect 39 556 40 558
rect 42 556 43 558
rect 31 465 35 466
rect 31 463 32 465
rect 34 463 35 465
rect 31 461 35 463
rect 31 459 32 461
rect 34 459 35 461
rect 31 458 35 459
rect 28 453 32 454
rect 28 451 29 453
rect 31 451 32 453
rect 28 415 32 451
rect 28 413 29 415
rect 31 413 32 415
rect 28 412 32 413
rect 39 270 43 556
rect 47 686 119 687
rect 47 684 116 686
rect 118 684 119 686
rect 47 683 119 684
rect 47 605 51 683
rect 55 678 87 679
rect 257 678 261 695
rect 324 695 328 708
rect 614 710 664 711
rect 614 708 661 710
rect 663 708 664 710
rect 614 707 664 708
rect 614 703 618 707
rect 614 701 615 703
rect 617 701 618 703
rect 614 700 618 701
rect 660 702 664 703
rect 660 700 661 702
rect 663 700 664 702
rect 324 693 325 695
rect 327 693 328 695
rect 324 692 328 693
rect 478 694 529 698
rect 289 685 332 686
rect 289 683 290 685
rect 292 683 332 685
rect 289 682 332 683
rect 55 676 84 678
rect 86 676 87 678
rect 55 675 87 676
rect 167 677 171 678
rect 167 675 168 677
rect 170 675 171 677
rect 55 623 59 675
rect 104 673 108 674
rect 104 671 105 673
rect 107 671 108 673
rect 55 621 56 623
rect 58 621 59 623
rect 55 620 59 621
rect 83 667 108 671
rect 83 615 87 667
rect 167 665 171 675
rect 257 674 291 678
rect 185 669 219 670
rect 185 667 186 669
rect 188 667 219 669
rect 185 666 219 667
rect 132 661 171 665
rect 95 644 99 645
rect 95 642 96 644
rect 98 642 99 644
rect 95 628 99 642
rect 95 626 96 628
rect 98 626 99 628
rect 95 624 99 626
rect 114 622 122 623
rect 114 620 115 622
rect 117 620 119 622
rect 121 620 122 622
rect 114 619 122 620
rect 83 613 84 615
rect 86 613 87 615
rect 83 611 87 613
rect 119 608 128 609
rect 119 606 120 608
rect 122 606 125 608
rect 127 606 128 608
rect 119 605 128 606
rect 47 603 48 605
rect 50 603 51 605
rect 47 402 51 603
rect 132 598 136 661
rect 152 644 211 645
rect 152 642 153 644
rect 155 642 211 644
rect 152 641 211 642
rect 207 638 211 641
rect 207 636 208 638
rect 210 636 211 638
rect 207 635 211 636
rect 148 630 205 631
rect 148 628 149 630
rect 151 628 205 630
rect 148 627 205 628
rect 215 630 219 666
rect 287 644 291 674
rect 287 642 288 644
rect 290 642 291 644
rect 287 641 291 642
rect 317 677 321 678
rect 317 675 318 677
rect 320 675 321 677
rect 215 628 216 630
rect 218 628 219 630
rect 215 627 219 628
rect 201 623 205 627
rect 171 622 175 623
rect 171 620 172 622
rect 174 620 175 622
rect 67 597 136 598
rect 67 595 68 597
rect 70 595 136 597
rect 67 594 136 595
rect 163 605 167 606
rect 163 603 164 605
rect 166 603 167 605
rect 107 574 111 594
rect 163 584 167 603
rect 163 582 164 584
rect 166 582 167 584
rect 163 581 167 582
rect 171 584 175 620
rect 201 622 227 623
rect 201 620 224 622
rect 226 620 227 622
rect 201 619 227 620
rect 180 608 184 609
rect 317 608 321 675
rect 180 606 181 608
rect 183 606 184 608
rect 271 607 321 608
rect 180 605 184 606
rect 180 603 181 605
rect 183 603 184 605
rect 180 592 184 603
rect 248 606 252 607
rect 248 604 249 606
rect 251 604 252 606
rect 271 605 272 607
rect 274 605 321 607
rect 271 604 321 605
rect 248 600 252 604
rect 248 599 299 600
rect 248 597 296 599
rect 298 597 299 599
rect 248 596 299 597
rect 180 591 291 592
rect 180 589 288 591
rect 290 589 291 591
rect 180 588 291 589
rect 171 582 172 584
rect 174 582 175 584
rect 171 581 175 582
rect 107 572 108 574
rect 110 572 111 574
rect 107 570 111 572
rect 154 566 259 567
rect 84 565 150 566
rect 84 563 85 565
rect 87 563 150 565
rect 154 564 155 566
rect 157 564 256 566
rect 258 564 259 566
rect 154 563 259 564
rect 84 562 150 563
rect 146 558 150 562
rect 328 559 332 682
rect 55 557 115 558
rect 55 555 88 557
rect 90 555 112 557
rect 114 555 115 557
rect 146 556 147 558
rect 149 556 150 558
rect 146 555 150 556
rect 223 558 332 559
rect 223 556 224 558
rect 226 556 332 558
rect 223 555 332 556
rect 55 554 115 555
rect 55 479 59 554
rect 240 550 324 551
rect 240 548 241 550
rect 243 548 321 550
rect 323 548 324 550
rect 240 547 324 548
rect 187 542 211 543
rect 55 477 56 479
rect 58 477 59 479
rect 55 476 59 477
rect 91 541 122 542
rect 91 539 119 541
rect 121 539 122 541
rect 187 540 188 542
rect 190 540 211 542
rect 187 539 211 540
rect 91 538 122 539
rect 91 472 95 538
rect 195 534 203 535
rect 99 533 103 534
rect 99 531 100 533
rect 102 531 103 533
rect 195 532 196 534
rect 198 532 203 534
rect 195 531 203 532
rect 99 500 103 531
rect 99 498 100 500
rect 102 498 103 500
rect 99 497 103 498
rect 199 494 203 531
rect 207 501 211 539
rect 222 534 226 535
rect 222 532 223 534
rect 225 532 226 534
rect 222 530 226 532
rect 222 528 223 530
rect 225 528 226 530
rect 222 527 226 528
rect 207 497 254 501
rect 199 492 200 494
rect 202 492 203 494
rect 199 490 203 492
rect 219 487 226 488
rect 99 486 131 487
rect 99 484 100 486
rect 102 484 128 486
rect 130 484 131 486
rect 219 485 220 487
rect 222 485 223 487
rect 225 485 226 487
rect 219 484 226 485
rect 99 483 131 484
rect 250 483 254 497
rect 259 487 315 488
rect 259 485 260 487
rect 262 485 315 487
rect 259 484 315 485
rect 250 481 251 483
rect 253 481 254 483
rect 250 480 254 481
rect 55 471 95 472
rect 55 469 56 471
rect 58 469 95 471
rect 55 468 95 469
rect 95 462 194 463
rect 55 461 79 462
rect 55 459 56 461
rect 58 459 72 461
rect 74 459 76 461
rect 78 459 79 461
rect 95 460 96 462
rect 98 460 191 462
rect 193 460 194 462
rect 95 459 194 460
rect 220 461 231 462
rect 220 459 221 461
rect 223 459 228 461
rect 230 459 231 461
rect 55 458 79 459
rect 220 458 231 459
rect 67 453 140 454
rect 67 451 68 453
rect 70 451 136 453
rect 138 451 140 453
rect 67 450 140 451
rect 71 438 299 439
rect 71 436 72 438
rect 74 436 296 438
rect 298 436 299 438
rect 71 435 299 436
rect 99 428 279 429
rect 99 426 100 428
rect 102 426 276 428
rect 278 426 279 428
rect 99 425 279 426
rect 107 420 111 421
rect 107 418 108 420
rect 110 418 111 420
rect 56 415 96 416
rect 56 413 57 415
rect 59 413 92 415
rect 94 413 96 415
rect 56 412 96 413
rect 47 400 48 402
rect 50 400 51 402
rect 47 399 51 400
rect 90 398 94 399
rect 90 396 91 398
rect 93 396 94 398
rect 90 394 94 396
rect 52 390 94 394
rect 52 346 56 390
rect 67 384 94 385
rect 67 382 68 384
rect 70 382 94 384
rect 67 381 94 382
rect 52 344 53 346
rect 55 344 56 346
rect 52 343 56 344
rect 63 376 67 377
rect 63 374 64 376
rect 66 374 67 376
rect 63 343 67 374
rect 63 341 64 343
rect 66 341 67 343
rect 63 340 67 341
rect 67 334 71 335
rect 67 332 68 334
rect 70 332 71 334
rect 39 268 40 270
rect 42 268 43 270
rect 39 145 43 268
rect 47 318 51 319
rect 47 316 48 318
rect 50 316 51 318
rect 47 314 51 316
rect 47 312 48 314
rect 50 312 51 314
rect 47 195 51 312
rect 67 309 71 332
rect 90 326 94 381
rect 107 341 111 418
rect 131 420 271 421
rect 131 418 132 420
rect 134 418 271 420
rect 131 417 271 418
rect 267 415 271 417
rect 267 413 268 415
rect 270 413 271 415
rect 140 412 175 413
rect 140 410 141 412
rect 143 410 172 412
rect 174 410 175 412
rect 140 409 175 410
rect 205 412 219 413
rect 267 412 271 413
rect 205 410 206 412
rect 208 410 216 412
rect 218 410 219 412
rect 205 409 219 410
rect 179 406 183 407
rect 179 404 180 406
rect 182 404 183 406
rect 107 339 108 341
rect 110 339 111 341
rect 107 338 111 339
rect 116 393 120 394
rect 116 391 117 393
rect 119 391 120 393
rect 90 324 91 326
rect 93 324 94 326
rect 90 323 94 324
rect 116 322 120 391
rect 162 390 173 391
rect 148 389 158 390
rect 148 387 149 389
rect 151 387 155 389
rect 157 387 158 389
rect 148 386 158 387
rect 162 388 170 390
rect 172 388 173 390
rect 162 387 173 388
rect 131 376 135 377
rect 131 374 132 376
rect 134 374 135 376
rect 131 343 135 374
rect 131 341 132 343
rect 134 341 135 343
rect 131 340 135 341
rect 148 356 152 357
rect 148 354 149 356
rect 151 354 152 356
rect 148 326 152 354
rect 162 340 166 387
rect 162 338 163 340
rect 165 338 166 340
rect 162 337 166 338
rect 179 340 183 404
rect 231 405 235 406
rect 231 403 232 405
rect 234 403 235 405
rect 231 402 235 403
rect 201 401 235 402
rect 201 399 202 401
rect 204 399 235 401
rect 201 398 235 399
rect 275 398 279 425
rect 275 396 276 398
rect 278 396 279 398
rect 275 395 279 396
rect 311 406 315 484
rect 311 404 312 406
rect 314 404 315 406
rect 243 393 247 394
rect 243 391 244 393
rect 246 391 247 393
rect 243 377 247 391
rect 288 382 292 383
rect 288 380 289 382
rect 291 380 292 382
rect 179 338 180 340
rect 182 338 183 340
rect 179 337 183 338
rect 220 376 224 377
rect 220 374 221 376
rect 223 374 224 376
rect 220 336 224 374
rect 243 373 271 377
rect 231 356 235 357
rect 231 354 232 356
rect 234 354 235 356
rect 231 343 235 354
rect 231 341 232 343
rect 234 341 235 343
rect 231 340 235 341
rect 211 335 230 336
rect 211 333 212 335
rect 214 333 227 335
rect 229 333 230 335
rect 211 332 230 333
rect 148 324 149 326
rect 151 324 152 326
rect 148 323 152 324
rect 267 326 271 373
rect 288 344 292 380
rect 284 343 292 344
rect 284 341 285 343
rect 287 341 292 343
rect 284 340 292 341
rect 267 324 268 326
rect 270 324 271 326
rect 267 323 271 324
rect 116 320 117 322
rect 119 320 120 322
rect 116 318 120 320
rect 204 317 208 318
rect 204 315 205 317
rect 207 315 208 317
rect 67 307 68 309
rect 70 307 71 309
rect 67 306 71 307
rect 75 309 79 310
rect 75 307 76 309
rect 78 307 79 309
rect 75 284 79 307
rect 204 305 208 315
rect 231 317 256 318
rect 231 315 232 317
rect 234 315 253 317
rect 255 315 256 317
rect 231 314 256 315
rect 311 305 315 404
rect 75 282 76 284
rect 78 282 79 284
rect 75 281 79 282
rect 166 301 315 305
rect 320 390 324 547
rect 320 388 321 390
rect 323 388 324 390
rect 87 278 148 279
rect 87 276 88 278
rect 90 276 148 278
rect 87 275 148 276
rect 144 262 148 275
rect 99 261 103 262
rect 99 259 100 261
rect 102 259 103 261
rect 144 260 145 262
rect 147 260 148 262
rect 144 259 148 260
rect 166 262 170 301
rect 213 284 283 285
rect 213 282 214 284
rect 216 282 283 284
rect 213 281 283 282
rect 191 270 217 271
rect 191 268 192 270
rect 194 268 214 270
rect 216 268 217 270
rect 191 267 217 268
rect 279 270 283 281
rect 279 268 280 270
rect 282 268 283 270
rect 279 267 283 268
rect 166 260 167 262
rect 169 260 170 262
rect 47 193 48 195
rect 50 193 51 195
rect 47 167 51 193
rect 64 246 86 247
rect 64 244 83 246
rect 85 244 86 246
rect 64 243 86 244
rect 64 191 68 243
rect 99 239 103 259
rect 166 255 170 260
rect 127 254 170 255
rect 127 252 128 254
rect 130 252 170 254
rect 127 251 170 252
rect 64 189 65 191
rect 67 189 68 191
rect 64 188 68 189
rect 75 235 103 239
rect 159 246 163 247
rect 159 244 160 246
rect 162 244 163 246
rect 75 175 79 235
rect 159 213 163 244
rect 279 246 316 248
rect 279 244 280 246
rect 282 244 316 246
rect 279 243 316 244
rect 97 209 163 213
rect 204 237 208 238
rect 204 235 205 237
rect 207 235 208 237
rect 97 194 101 209
rect 108 198 169 199
rect 108 196 109 198
rect 111 196 169 198
rect 204 197 208 235
rect 108 195 169 196
rect 97 192 98 194
rect 100 192 101 194
rect 97 191 101 192
rect 143 190 147 191
rect 143 188 144 190
rect 146 188 147 190
rect 56 174 79 175
rect 56 172 57 174
rect 59 172 79 174
rect 56 171 79 172
rect 83 182 87 183
rect 83 180 84 182
rect 86 180 87 182
rect 83 167 87 180
rect 47 163 87 167
rect 135 174 139 175
rect 135 172 136 174
rect 138 172 139 174
rect 135 160 139 172
rect 135 158 136 160
rect 138 158 139 160
rect 135 157 139 158
rect 143 161 147 188
rect 165 174 169 195
rect 173 196 208 197
rect 173 194 174 196
rect 176 194 208 196
rect 173 193 208 194
rect 226 220 230 221
rect 226 218 227 220
rect 229 218 230 220
rect 226 183 230 218
rect 165 172 166 174
rect 168 172 169 174
rect 165 171 169 172
rect 215 182 230 183
rect 215 180 216 182
rect 218 180 230 182
rect 215 179 230 180
rect 143 160 201 161
rect 143 158 198 160
rect 200 158 201 160
rect 143 157 201 158
rect 39 144 211 145
rect 39 142 208 144
rect 210 142 211 144
rect 39 141 211 142
rect 39 127 43 141
rect 99 135 148 136
rect 99 133 100 135
rect 102 133 136 135
rect 138 133 148 135
rect 99 132 148 133
rect 144 127 148 132
rect 39 125 40 127
rect 42 125 43 127
rect 39 124 43 125
rect 87 126 111 127
rect 87 124 88 126
rect 90 124 108 126
rect 110 124 111 126
rect 144 125 145 127
rect 147 125 148 127
rect 144 124 148 125
rect 87 123 111 124
rect 197 119 201 120
rect 197 117 198 119
rect 200 117 201 119
rect 197 114 201 117
rect 150 112 173 113
rect 150 110 170 112
rect 172 110 173 112
rect 116 109 120 110
rect 116 107 117 109
rect 119 107 120 109
rect 41 101 84 102
rect 41 99 81 101
rect 83 99 84 101
rect 41 98 84 99
rect 31 88 35 89
rect 31 86 32 88
rect 34 86 35 88
rect 31 46 35 86
rect 31 44 32 46
rect 34 44 35 46
rect 31 43 35 44
rect 41 30 45 98
rect 116 94 120 107
rect 150 109 173 110
rect 197 112 198 114
rect 200 112 201 114
rect 64 90 120 94
rect 137 101 141 102
rect 137 99 138 101
rect 140 99 141 101
rect 64 47 68 90
rect 137 54 141 99
rect 89 53 141 54
rect 89 51 90 53
rect 92 51 141 53
rect 89 50 141 51
rect 64 45 65 47
rect 67 45 68 47
rect 64 44 68 45
rect 150 39 154 109
rect 189 102 193 104
rect 189 100 190 102
rect 192 100 193 102
rect 189 64 193 100
rect 166 63 193 64
rect 166 61 167 63
rect 169 61 193 63
rect 166 60 193 61
rect 197 54 201 112
rect 197 52 198 54
rect 200 52 201 54
rect 197 51 201 52
rect 207 47 211 141
rect 215 88 219 179
rect 312 153 316 243
rect 320 169 324 388
rect 320 167 321 169
rect 323 167 324 169
rect 320 166 324 167
rect 328 415 332 555
rect 328 413 329 415
rect 331 413 332 415
rect 328 160 332 413
rect 328 158 329 160
rect 331 158 332 160
rect 328 157 332 158
rect 355 577 438 581
rect 355 153 360 577
rect 312 149 360 153
rect 347 148 360 149
rect 373 572 377 573
rect 373 570 374 572
rect 376 570 377 572
rect 373 317 377 570
rect 373 315 374 317
rect 376 315 377 317
rect 373 175 377 315
rect 381 563 385 564
rect 381 561 382 563
rect 384 561 385 563
rect 381 342 385 561
rect 434 552 438 577
rect 478 568 482 694
rect 525 687 529 694
rect 521 686 529 687
rect 521 684 522 686
rect 524 684 529 686
rect 521 683 529 684
rect 551 693 555 694
rect 551 691 552 693
rect 554 691 555 693
rect 504 678 508 679
rect 504 676 505 678
rect 507 676 508 678
rect 442 567 482 568
rect 442 565 443 567
rect 445 565 482 567
rect 442 564 482 565
rect 486 644 490 645
rect 486 642 487 644
rect 489 642 490 644
rect 434 551 462 552
rect 486 551 490 642
rect 504 618 508 676
rect 512 669 539 670
rect 512 667 536 669
rect 538 667 539 669
rect 512 666 539 667
rect 512 630 516 666
rect 512 628 513 630
rect 515 628 516 630
rect 512 626 516 628
rect 551 621 555 691
rect 637 685 641 686
rect 637 683 638 685
rect 640 683 641 685
rect 564 679 616 680
rect 564 677 613 679
rect 615 677 616 679
rect 564 676 616 677
rect 564 631 568 676
rect 637 640 641 683
rect 564 629 565 631
rect 567 629 568 631
rect 564 628 568 629
rect 585 636 641 640
rect 504 616 505 618
rect 507 616 508 618
rect 532 620 555 621
rect 585 623 589 636
rect 660 632 664 700
rect 670 686 674 687
rect 670 684 671 686
rect 673 684 674 686
rect 670 644 674 684
rect 670 642 671 644
rect 673 642 674 644
rect 670 641 674 642
rect 621 631 664 632
rect 621 629 622 631
rect 624 629 664 631
rect 621 628 664 629
rect 585 621 586 623
rect 588 621 589 623
rect 585 620 589 621
rect 532 618 533 620
rect 535 618 555 620
rect 532 617 555 618
rect 504 613 508 616
rect 504 611 505 613
rect 507 611 508 613
rect 504 610 508 611
rect 594 606 618 607
rect 557 605 561 606
rect 557 603 558 605
rect 560 603 561 605
rect 594 604 595 606
rect 597 604 615 606
rect 617 604 618 606
rect 594 603 618 604
rect 662 605 666 606
rect 662 603 663 605
rect 665 603 666 605
rect 557 598 561 603
rect 557 597 606 598
rect 557 595 567 597
rect 569 595 603 597
rect 605 595 606 597
rect 557 594 606 595
rect 662 589 666 603
rect 494 588 666 589
rect 494 586 495 588
rect 497 586 666 588
rect 494 585 666 586
rect 504 572 562 573
rect 504 570 505 572
rect 507 570 562 572
rect 504 569 562 570
rect 434 549 459 551
rect 461 549 462 551
rect 434 548 462 549
rect 475 550 490 551
rect 475 548 487 550
rect 489 548 490 550
rect 475 547 490 548
rect 536 558 540 559
rect 536 556 537 558
rect 539 556 540 558
rect 475 512 479 547
rect 475 510 476 512
rect 478 510 479 512
rect 475 509 479 510
rect 497 536 532 537
rect 497 534 529 536
rect 531 534 532 536
rect 497 533 532 534
rect 536 535 540 556
rect 558 542 562 569
rect 566 572 570 573
rect 566 570 567 572
rect 569 570 570 572
rect 566 558 570 570
rect 566 556 567 558
rect 569 556 570 558
rect 566 555 570 556
rect 618 563 658 567
rect 618 550 622 563
rect 618 548 619 550
rect 621 548 622 550
rect 618 547 622 548
rect 626 558 649 559
rect 626 556 646 558
rect 648 556 649 558
rect 626 555 649 556
rect 558 540 559 542
rect 561 540 562 542
rect 558 539 562 540
rect 604 538 608 539
rect 604 536 605 538
rect 607 536 608 538
rect 536 534 597 535
rect 497 495 501 533
rect 536 532 594 534
rect 596 532 597 534
rect 536 531 597 532
rect 604 521 608 536
rect 497 493 498 495
rect 500 493 501 495
rect 497 492 501 493
rect 542 517 608 521
rect 542 486 546 517
rect 626 495 630 555
rect 542 484 543 486
rect 545 484 546 486
rect 542 483 546 484
rect 602 491 630 495
rect 637 541 641 542
rect 637 539 638 541
rect 640 539 641 541
rect 535 478 578 479
rect 535 476 575 478
rect 577 476 578 478
rect 535 475 578 476
rect 535 470 539 475
rect 602 471 606 491
rect 637 487 641 539
rect 619 486 641 487
rect 619 484 620 486
rect 622 484 641 486
rect 619 483 641 484
rect 654 537 658 563
rect 654 535 655 537
rect 657 535 658 537
rect 535 468 536 470
rect 538 468 539 470
rect 488 462 514 463
rect 488 460 489 462
rect 491 460 511 462
rect 513 460 514 462
rect 488 459 514 460
rect 535 429 539 468
rect 557 470 561 471
rect 557 468 558 470
rect 560 468 561 470
rect 602 469 603 471
rect 605 469 606 471
rect 602 468 606 469
rect 557 455 561 468
rect 557 454 618 455
rect 557 452 615 454
rect 617 452 618 454
rect 557 451 618 452
rect 381 340 382 342
rect 384 340 385 342
rect 381 183 385 340
rect 390 425 539 429
rect 390 326 394 425
rect 449 415 474 416
rect 449 413 450 415
rect 452 413 471 415
rect 473 413 474 415
rect 449 412 474 413
rect 497 415 501 425
rect 497 413 498 415
rect 500 413 501 415
rect 497 412 501 413
rect 634 423 638 424
rect 634 421 635 423
rect 637 421 638 423
rect 585 410 589 412
rect 585 408 586 410
rect 588 408 589 410
rect 434 406 438 407
rect 434 404 435 406
rect 437 404 438 406
rect 413 389 421 390
rect 413 387 418 389
rect 420 387 421 389
rect 413 386 421 387
rect 413 350 417 386
rect 434 357 438 404
rect 553 406 557 407
rect 553 404 554 406
rect 556 404 557 406
rect 475 397 494 398
rect 475 395 476 397
rect 478 395 491 397
rect 493 395 494 397
rect 475 394 494 395
rect 470 389 474 390
rect 470 387 471 389
rect 473 387 474 389
rect 470 376 474 387
rect 470 374 471 376
rect 473 374 474 376
rect 470 373 474 374
rect 434 353 462 357
rect 481 356 485 394
rect 481 354 482 356
rect 484 354 485 356
rect 481 353 485 354
rect 522 392 526 393
rect 522 390 523 392
rect 525 390 526 392
rect 413 348 414 350
rect 416 348 417 350
rect 413 347 417 348
rect 458 339 462 353
rect 458 337 459 339
rect 461 337 462 339
rect 458 336 462 337
rect 390 324 391 326
rect 393 324 394 326
rect 390 246 394 324
rect 426 334 430 335
rect 426 332 427 334
rect 429 332 430 334
rect 426 305 430 332
rect 470 331 504 332
rect 470 329 501 331
rect 503 329 504 331
rect 470 328 504 329
rect 470 327 474 328
rect 470 325 471 327
rect 473 325 474 327
rect 470 324 474 325
rect 522 326 526 390
rect 539 392 543 393
rect 539 390 540 392
rect 542 390 543 392
rect 539 343 543 390
rect 553 376 557 404
rect 553 374 554 376
rect 556 374 557 376
rect 553 373 557 374
rect 570 389 574 390
rect 570 387 571 389
rect 573 387 574 389
rect 570 356 574 387
rect 570 354 571 356
rect 573 354 574 356
rect 570 353 574 354
rect 532 342 543 343
rect 532 340 533 342
rect 535 340 543 342
rect 547 343 557 344
rect 547 341 548 343
rect 550 341 554 343
rect 556 341 557 343
rect 547 340 557 341
rect 532 339 543 340
rect 585 339 589 408
rect 611 406 615 407
rect 611 404 612 406
rect 614 404 615 406
rect 585 337 586 339
rect 588 337 589 339
rect 585 336 589 337
rect 594 391 598 392
rect 594 389 595 391
rect 597 389 598 391
rect 522 324 523 326
rect 525 324 526 326
rect 522 323 526 324
rect 486 320 500 321
rect 486 318 487 320
rect 489 318 497 320
rect 499 318 500 320
rect 434 317 438 318
rect 486 317 500 318
rect 530 320 565 321
rect 530 318 531 320
rect 533 318 562 320
rect 564 318 565 320
rect 530 317 565 318
rect 434 315 435 317
rect 437 315 438 317
rect 434 313 438 315
rect 434 312 574 313
rect 434 310 571 312
rect 573 310 574 312
rect 434 309 574 310
rect 594 312 598 389
rect 611 349 615 404
rect 634 398 638 421
rect 654 418 658 535
rect 654 416 655 418
rect 657 416 658 418
rect 654 414 658 416
rect 654 412 655 414
rect 657 412 658 414
rect 654 411 658 412
rect 662 462 666 585
rect 662 460 663 462
rect 665 460 666 462
rect 634 396 635 398
rect 637 396 638 398
rect 634 395 638 396
rect 638 389 642 390
rect 638 387 639 389
rect 641 387 642 389
rect 638 356 642 387
rect 638 354 639 356
rect 641 354 642 356
rect 638 353 642 354
rect 649 386 653 387
rect 649 384 650 386
rect 652 384 653 386
rect 611 348 638 349
rect 611 346 635 348
rect 637 346 638 348
rect 611 345 638 346
rect 649 340 653 384
rect 611 336 653 340
rect 611 334 615 336
rect 611 332 612 334
rect 614 332 615 334
rect 611 331 615 332
rect 654 330 658 331
rect 654 328 655 330
rect 657 328 658 330
rect 609 317 649 318
rect 609 315 611 317
rect 613 315 646 317
rect 648 315 649 317
rect 609 314 649 315
rect 594 310 595 312
rect 597 310 598 312
rect 594 309 598 310
rect 426 304 606 305
rect 426 302 427 304
rect 429 302 603 304
rect 605 302 606 304
rect 426 301 606 302
rect 406 294 634 295
rect 406 292 407 294
rect 409 292 631 294
rect 633 292 634 294
rect 406 291 634 292
rect 565 279 638 280
rect 565 277 567 279
rect 569 277 635 279
rect 637 277 638 279
rect 565 276 638 277
rect 474 271 485 272
rect 626 271 650 272
rect 474 269 475 271
rect 477 269 482 271
rect 484 269 485 271
rect 474 268 485 269
rect 511 270 610 271
rect 511 268 512 270
rect 514 268 607 270
rect 609 268 610 270
rect 626 269 627 271
rect 629 269 631 271
rect 633 269 647 271
rect 649 269 650 271
rect 626 268 650 269
rect 511 267 610 268
rect 610 261 650 262
rect 610 259 647 261
rect 649 259 650 261
rect 610 258 650 259
rect 451 249 455 250
rect 451 247 452 249
rect 454 247 455 249
rect 390 245 446 246
rect 390 243 443 245
rect 445 243 446 245
rect 390 242 446 243
rect 451 233 455 247
rect 574 246 606 247
rect 479 245 486 246
rect 479 243 480 245
rect 482 243 483 245
rect 485 243 486 245
rect 574 244 575 246
rect 577 244 603 246
rect 605 244 606 246
rect 574 243 606 244
rect 479 242 486 243
rect 502 238 506 240
rect 502 236 503 238
rect 505 236 506 238
rect 451 229 498 233
rect 479 202 483 203
rect 479 200 480 202
rect 482 200 483 202
rect 479 198 483 200
rect 479 196 480 198
rect 482 196 483 198
rect 479 195 483 196
rect 494 191 498 229
rect 502 199 506 236
rect 602 232 606 233
rect 602 230 603 232
rect 605 230 606 232
rect 602 199 606 230
rect 502 198 510 199
rect 502 196 507 198
rect 509 196 510 198
rect 602 197 603 199
rect 605 197 606 199
rect 602 196 606 197
rect 502 195 510 196
rect 610 192 614 258
rect 583 191 614 192
rect 494 190 518 191
rect 494 188 515 190
rect 517 188 518 190
rect 583 189 584 191
rect 586 189 614 191
rect 583 188 614 189
rect 646 253 650 254
rect 646 251 647 253
rect 649 251 650 253
rect 494 187 518 188
rect 381 182 465 183
rect 381 180 382 182
rect 384 180 462 182
rect 464 180 465 182
rect 381 179 465 180
rect 646 176 650 251
rect 590 175 650 176
rect 373 174 482 175
rect 373 172 479 174
rect 481 172 482 174
rect 373 171 482 172
rect 555 174 559 175
rect 555 172 556 174
rect 558 172 559 174
rect 590 173 591 175
rect 593 173 615 175
rect 617 173 650 175
rect 590 172 650 173
rect 215 86 216 88
rect 218 86 219 88
rect 215 85 219 86
rect 189 46 211 47
rect 189 44 190 46
rect 192 44 211 46
rect 373 48 377 171
rect 555 168 559 172
rect 555 167 621 168
rect 446 166 551 167
rect 446 164 447 166
rect 449 164 548 166
rect 550 164 551 166
rect 555 165 618 167
rect 620 165 621 167
rect 555 164 621 165
rect 446 163 551 164
rect 594 158 598 160
rect 594 156 595 158
rect 597 156 598 158
rect 530 148 534 149
rect 530 146 531 148
rect 533 146 534 148
rect 414 141 525 142
rect 414 139 415 141
rect 417 139 525 141
rect 414 138 525 139
rect 406 133 457 134
rect 406 131 407 133
rect 409 131 457 133
rect 406 130 457 131
rect 453 126 457 130
rect 384 125 434 126
rect 384 123 431 125
rect 433 123 434 125
rect 453 124 454 126
rect 456 124 457 126
rect 453 123 457 124
rect 521 127 525 138
rect 521 125 522 127
rect 524 125 525 127
rect 521 124 525 125
rect 384 122 434 123
rect 521 122 522 124
rect 524 122 525 124
rect 384 55 388 122
rect 521 121 525 122
rect 478 110 504 111
rect 478 108 479 110
rect 481 108 504 110
rect 478 107 504 108
rect 530 110 534 146
rect 538 148 542 149
rect 538 146 539 148
rect 541 146 542 148
rect 538 127 542 146
rect 594 136 598 156
rect 538 125 539 127
rect 541 125 542 127
rect 538 124 542 125
rect 569 135 638 136
rect 569 133 635 135
rect 637 133 638 135
rect 569 132 638 133
rect 530 108 531 110
rect 533 108 534 110
rect 530 107 534 108
rect 500 103 504 107
rect 486 102 490 103
rect 486 100 487 102
rect 489 100 490 102
rect 384 53 385 55
rect 387 53 388 55
rect 384 52 388 53
rect 414 88 418 89
rect 414 86 415 88
rect 417 86 418 88
rect 414 56 418 86
rect 486 64 490 100
rect 500 102 557 103
rect 500 100 554 102
rect 556 100 557 102
rect 500 99 557 100
rect 494 94 498 95
rect 494 92 495 94
rect 497 92 498 94
rect 494 89 498 92
rect 494 88 553 89
rect 494 86 550 88
rect 552 86 553 88
rect 494 85 553 86
rect 569 69 573 132
rect 654 127 658 328
rect 654 125 655 127
rect 657 125 658 127
rect 577 124 586 125
rect 577 122 578 124
rect 580 122 583 124
rect 585 122 586 124
rect 577 121 586 122
rect 618 117 622 119
rect 618 115 619 117
rect 621 115 622 117
rect 583 110 591 111
rect 583 108 584 110
rect 586 108 588 110
rect 590 108 591 110
rect 583 107 591 108
rect 606 104 610 106
rect 606 102 607 104
rect 609 102 610 104
rect 606 88 610 102
rect 606 86 607 88
rect 609 86 610 88
rect 606 85 610 86
rect 534 65 573 69
rect 486 63 520 64
rect 486 61 517 63
rect 519 61 520 63
rect 486 60 520 61
rect 414 52 448 56
rect 534 55 538 65
rect 618 63 622 115
rect 597 59 622 63
rect 646 109 650 110
rect 646 107 647 109
rect 649 107 650 109
rect 597 57 598 59
rect 600 57 601 59
rect 597 56 601 57
rect 646 55 650 107
rect 534 53 535 55
rect 537 53 538 55
rect 534 52 538 53
rect 618 54 650 55
rect 618 52 619 54
rect 621 52 650 54
rect 373 47 416 48
rect 373 45 413 47
rect 415 45 416 47
rect 373 44 416 45
rect 189 43 211 44
rect 150 37 151 39
rect 153 37 154 39
rect 150 36 154 37
rect 377 37 381 38
rect 377 35 378 37
rect 380 35 381 37
rect 41 28 42 30
rect 44 28 45 30
rect 41 27 45 28
rect 87 29 91 30
rect 87 27 88 29
rect 90 27 91 29
rect 87 23 91 27
rect 41 22 91 23
rect 41 20 42 22
rect 44 20 91 22
rect 41 19 91 20
rect 377 22 381 35
rect 444 35 448 52
rect 618 51 650 52
rect 654 47 658 125
rect 586 46 658 47
rect 586 44 587 46
rect 589 44 658 46
rect 586 43 658 44
rect 662 174 666 460
rect 673 317 677 318
rect 673 315 674 317
rect 676 315 677 317
rect 673 279 677 315
rect 673 277 674 279
rect 676 277 677 279
rect 673 276 677 277
rect 670 271 674 272
rect 670 269 671 271
rect 673 269 674 271
rect 670 267 674 269
rect 670 265 671 267
rect 673 265 674 267
rect 670 264 674 265
rect 662 172 663 174
rect 665 172 666 174
rect 444 33 445 35
rect 447 33 448 35
rect 403 32 416 33
rect 444 32 448 33
rect 541 36 545 37
rect 541 34 542 36
rect 544 34 545 36
rect 541 32 545 34
rect 403 30 404 32
rect 406 30 413 32
rect 415 30 416 32
rect 541 30 542 32
rect 544 30 545 32
rect 662 30 666 172
rect 670 140 674 141
rect 670 138 671 140
rect 673 138 674 140
rect 670 125 674 138
rect 670 123 671 125
rect 673 123 674 125
rect 670 122 674 123
rect 403 29 416 30
rect 428 29 440 30
rect 428 27 429 29
rect 431 27 437 29
rect 439 27 440 29
rect 428 26 440 27
rect 514 29 518 30
rect 541 29 545 30
rect 586 29 618 30
rect 514 27 515 29
rect 517 27 518 29
rect 514 24 518 27
rect 586 27 587 29
rect 589 27 615 29
rect 617 27 618 29
rect 586 26 618 27
rect 662 28 663 30
rect 665 28 666 30
rect 662 26 666 28
rect 514 23 562 24
rect 377 21 456 22
rect 377 19 453 21
rect 455 19 456 21
rect 514 21 559 23
rect 561 21 562 23
rect 514 20 562 21
rect 377 18 456 19
<< alu3 >>
rect 259 703 269 704
rect 259 701 266 703
rect 268 701 269 703
rect 259 700 269 701
rect 298 700 324 701
rect 160 696 164 697
rect 160 694 161 696
rect 163 694 164 696
rect 160 649 164 694
rect 160 645 193 649
rect 95 644 156 645
rect 95 642 96 644
rect 98 642 153 644
rect 155 642 156 644
rect 95 641 156 642
rect 23 622 118 623
rect 23 620 115 622
rect 117 620 118 622
rect 23 619 118 620
rect 23 366 27 619
rect 124 608 184 609
rect 124 606 125 608
rect 127 606 181 608
rect 183 606 184 608
rect 124 605 184 606
rect 189 593 193 645
rect 31 592 193 593
rect 31 590 32 592
rect 34 590 193 592
rect 31 589 193 590
rect 31 465 35 466
rect 31 463 32 465
rect 34 463 35 465
rect 31 462 35 463
rect 31 461 59 462
rect 31 459 56 461
rect 58 459 59 461
rect 31 458 59 459
rect 63 376 67 589
rect 107 574 111 575
rect 107 572 108 574
rect 110 572 111 574
rect 84 565 88 566
rect 84 563 85 565
rect 87 563 88 565
rect 71 461 75 462
rect 71 459 72 461
rect 74 459 75 461
rect 71 438 75 459
rect 71 436 72 438
rect 74 436 75 438
rect 71 435 75 436
rect 63 374 64 376
rect 66 374 67 376
rect 63 373 67 374
rect 84 366 88 563
rect 23 362 88 366
rect 99 500 103 501
rect 99 498 100 500
rect 102 498 103 500
rect 99 486 103 498
rect 99 484 100 486
rect 102 484 103 486
rect 99 428 103 484
rect 99 426 100 428
rect 102 426 103 428
rect 23 315 27 362
rect 99 357 103 426
rect 107 420 111 572
rect 107 418 108 420
rect 110 418 111 420
rect 107 417 111 418
rect 131 420 135 589
rect 259 585 263 700
rect 298 698 299 700
rect 301 698 324 700
rect 298 697 324 698
rect 163 584 167 585
rect 163 582 164 584
rect 166 582 167 584
rect 163 462 167 582
rect 171 584 263 585
rect 171 582 172 584
rect 174 582 263 584
rect 171 581 263 582
rect 222 530 226 531
rect 222 528 223 530
rect 225 528 226 530
rect 222 488 226 528
rect 259 488 263 581
rect 222 487 263 488
rect 222 485 223 487
rect 225 485 260 487
rect 262 485 263 487
rect 222 484 263 485
rect 287 644 291 645
rect 287 642 288 644
rect 290 642 291 644
rect 287 591 291 642
rect 287 589 288 591
rect 290 589 291 591
rect 163 461 224 462
rect 163 459 221 461
rect 223 459 224 461
rect 163 458 224 459
rect 131 418 132 420
rect 134 418 135 420
rect 131 376 135 418
rect 171 412 209 413
rect 171 410 172 412
rect 174 410 206 412
rect 208 410 209 412
rect 171 409 209 410
rect 154 389 161 390
rect 154 387 155 389
rect 157 387 161 389
rect 154 386 161 387
rect 131 374 132 376
rect 134 374 135 376
rect 131 373 135 374
rect 157 357 161 386
rect 220 376 224 458
rect 287 429 291 589
rect 295 599 299 600
rect 295 597 296 599
rect 298 597 299 599
rect 295 438 299 597
rect 320 550 324 697
rect 486 644 674 645
rect 486 642 487 644
rect 489 642 671 644
rect 673 642 674 644
rect 486 641 674 642
rect 504 618 508 619
rect 504 616 505 618
rect 507 616 508 618
rect 320 548 321 550
rect 323 548 324 550
rect 320 547 324 548
rect 347 588 498 589
rect 347 586 495 588
rect 497 586 498 588
rect 347 585 498 586
rect 295 436 296 438
rect 298 436 299 438
rect 295 435 299 436
rect 275 428 291 429
rect 275 426 276 428
rect 278 426 291 428
rect 275 425 291 426
rect 220 374 221 376
rect 223 374 224 376
rect 220 373 224 374
rect 67 356 152 357
rect 67 354 149 356
rect 151 354 152 356
rect 67 353 152 354
rect 157 356 235 357
rect 157 354 232 356
rect 234 354 235 356
rect 157 353 235 354
rect 67 334 71 353
rect 67 332 68 334
rect 70 332 71 334
rect 67 331 71 332
rect 226 335 230 336
rect 226 333 227 335
rect 229 333 230 335
rect 23 314 51 315
rect 23 312 48 314
rect 50 312 51 314
rect 23 311 51 312
rect 75 284 217 285
rect 75 282 76 284
rect 78 282 214 284
rect 216 282 217 284
rect 75 281 217 282
rect 226 220 230 333
rect 226 218 227 220
rect 229 218 230 220
rect 226 217 230 218
rect 135 169 324 170
rect 135 167 321 169
rect 323 167 324 169
rect 135 166 324 167
rect 135 160 139 166
rect 135 158 136 160
rect 138 158 139 160
rect 135 135 139 158
rect 135 133 136 135
rect 138 133 139 135
rect 135 132 139 133
rect 197 160 332 161
rect 197 158 198 160
rect 200 158 329 160
rect 331 158 332 160
rect 197 157 332 158
rect 197 114 201 157
rect 347 145 352 585
rect 504 573 508 616
rect 373 572 508 573
rect 373 570 374 572
rect 376 570 505 572
rect 507 570 508 572
rect 373 569 508 570
rect 566 597 570 598
rect 566 595 567 597
rect 569 595 570 597
rect 566 572 570 595
rect 566 570 567 572
rect 569 570 570 572
rect 566 564 570 570
rect 381 563 570 564
rect 381 561 382 563
rect 384 561 570 563
rect 381 560 570 561
rect 475 512 479 513
rect 475 510 476 512
rect 478 510 479 512
rect 475 397 479 510
rect 654 418 682 419
rect 654 416 655 418
rect 657 416 682 418
rect 654 415 682 416
rect 475 395 476 397
rect 478 395 479 397
rect 475 394 479 395
rect 634 398 638 399
rect 634 396 635 398
rect 637 396 638 398
rect 634 377 638 396
rect 470 376 548 377
rect 470 374 471 376
rect 473 374 548 376
rect 470 373 548 374
rect 553 376 638 377
rect 553 374 554 376
rect 556 374 638 376
rect 553 373 638 374
rect 481 356 485 357
rect 481 354 482 356
rect 484 354 485 356
rect 414 304 430 305
rect 414 302 427 304
rect 429 302 430 304
rect 414 301 430 302
rect 406 294 410 295
rect 406 292 407 294
rect 409 292 410 294
rect 207 144 352 145
rect 207 142 208 144
rect 210 142 352 144
rect 207 141 352 142
rect 381 182 385 183
rect 381 180 382 182
rect 384 180 385 182
rect 197 112 198 114
rect 200 112 201 114
rect 197 111 201 112
rect 31 88 219 89
rect 31 86 32 88
rect 34 86 216 88
rect 218 86 219 88
rect 31 85 219 86
rect 381 33 385 180
rect 406 133 410 292
rect 406 131 407 133
rect 409 131 410 133
rect 406 130 410 131
rect 414 141 418 301
rect 481 272 485 354
rect 544 344 548 373
rect 570 356 574 357
rect 570 354 571 356
rect 573 354 574 356
rect 544 343 551 344
rect 544 341 548 343
rect 550 341 551 343
rect 544 340 551 341
rect 496 320 534 321
rect 496 318 497 320
rect 499 318 531 320
rect 533 318 534 320
rect 496 317 534 318
rect 570 312 574 354
rect 570 310 571 312
rect 573 310 574 312
rect 481 271 542 272
rect 481 269 482 271
rect 484 269 542 271
rect 481 268 542 269
rect 414 139 415 141
rect 417 139 418 141
rect 414 88 418 139
rect 414 86 415 88
rect 417 86 418 88
rect 414 85 418 86
rect 442 245 483 246
rect 442 243 443 245
rect 445 243 480 245
rect 482 243 483 245
rect 442 242 483 243
rect 442 149 446 242
rect 479 202 483 242
rect 479 200 480 202
rect 482 200 483 202
rect 479 199 483 200
rect 442 148 534 149
rect 442 146 531 148
rect 533 146 534 148
rect 442 145 534 146
rect 538 148 542 268
rect 538 146 539 148
rect 541 146 542 148
rect 538 145 542 146
rect 381 32 407 33
rect 381 30 404 32
rect 406 30 407 32
rect 442 30 446 145
rect 570 141 574 310
rect 594 312 598 313
rect 594 310 595 312
rect 597 310 598 312
rect 594 158 598 310
rect 602 304 606 373
rect 678 368 682 415
rect 602 302 603 304
rect 605 302 606 304
rect 602 246 606 302
rect 602 244 603 246
rect 605 244 606 246
rect 602 232 606 244
rect 602 230 603 232
rect 605 230 606 232
rect 602 229 606 230
rect 617 364 682 368
rect 617 167 621 364
rect 638 356 642 357
rect 638 354 639 356
rect 641 354 642 356
rect 630 294 634 295
rect 630 292 631 294
rect 633 292 634 294
rect 630 271 634 292
rect 630 269 631 271
rect 633 269 634 271
rect 630 268 634 269
rect 617 165 618 167
rect 620 165 621 167
rect 617 164 621 165
rect 594 156 595 158
rect 597 156 598 158
rect 594 155 598 156
rect 638 141 642 354
rect 646 271 674 272
rect 646 269 647 271
rect 649 269 674 271
rect 646 268 674 269
rect 670 267 674 268
rect 670 265 671 267
rect 673 265 674 267
rect 670 264 674 265
rect 512 140 674 141
rect 512 138 671 140
rect 673 138 674 140
rect 512 137 674 138
rect 512 85 516 137
rect 521 124 581 125
rect 521 122 522 124
rect 524 122 578 124
rect 580 122 581 124
rect 521 121 581 122
rect 678 111 682 364
rect 587 110 682 111
rect 587 108 588 110
rect 590 108 682 110
rect 587 107 682 108
rect 549 88 610 89
rect 549 86 550 88
rect 552 86 607 88
rect 609 86 610 88
rect 549 85 610 86
rect 512 81 545 85
rect 541 36 545 81
rect 541 34 542 36
rect 544 34 545 36
rect 541 33 545 34
rect 381 29 407 30
rect 436 29 446 30
rect 436 27 437 29
rect 439 27 446 29
rect 436 26 446 27
<< ptie >>
rect 32 720 38 722
rect 32 718 34 720
rect 36 718 38 720
rect 32 716 38 718
rect 120 720 126 722
rect 120 718 122 720
rect 124 718 126 720
rect 120 716 126 718
rect 136 720 142 722
rect 136 718 138 720
rect 140 718 142 720
rect 136 716 142 718
rect 180 720 186 722
rect 180 718 182 720
rect 184 718 186 720
rect 180 716 186 718
rect 310 720 328 722
rect 310 718 312 720
rect 314 718 324 720
rect 326 718 328 720
rect 310 716 328 718
rect 498 720 524 722
rect 498 718 500 720
rect 502 718 520 720
rect 522 718 524 720
rect 498 716 524 718
rect 536 720 542 722
rect 536 718 538 720
rect 540 718 542 720
rect 536 716 542 718
rect 607 720 625 722
rect 607 718 609 720
rect 611 718 621 720
rect 623 718 625 720
rect 607 716 625 718
rect 631 720 637 722
rect 631 718 633 720
rect 635 718 637 720
rect 631 707 637 718
rect 68 588 86 590
rect 68 586 70 588
rect 72 586 82 588
rect 84 586 86 588
rect 68 584 86 586
rect 96 588 102 590
rect 96 586 98 588
rect 100 586 102 588
rect 96 584 102 586
rect 140 588 146 590
rect 140 586 142 588
rect 144 586 146 588
rect 140 584 146 586
rect 272 588 278 605
rect 272 586 274 588
rect 276 586 278 588
rect 272 584 278 586
rect 501 588 519 590
rect 501 586 503 588
rect 505 586 515 588
rect 517 586 519 588
rect 501 584 519 586
rect 533 588 539 590
rect 533 586 535 588
rect 537 586 539 588
rect 533 584 539 586
rect 667 588 673 590
rect 667 586 669 588
rect 671 586 673 588
rect 667 584 673 586
rect 32 576 38 578
rect 32 574 34 576
rect 36 574 38 576
rect 32 572 38 574
rect 144 576 150 578
rect 144 574 146 576
rect 148 574 150 576
rect 144 557 150 574
rect 252 576 258 578
rect 252 574 254 576
rect 256 574 258 576
rect 252 572 258 574
rect 443 576 461 578
rect 443 574 445 576
rect 447 574 457 576
rect 459 574 461 576
rect 443 572 461 574
rect 507 576 513 578
rect 507 574 509 576
rect 511 574 513 576
rect 507 563 513 574
rect 587 576 593 578
rect 587 574 589 576
rect 591 574 593 576
rect 587 572 593 574
rect 605 576 623 578
rect 605 574 607 576
rect 609 574 619 576
rect 621 574 623 576
rect 605 572 623 574
rect 631 576 637 578
rect 631 574 633 576
rect 635 574 637 576
rect 631 563 637 574
rect 52 444 58 446
rect 52 442 54 444
rect 56 442 58 444
rect 52 440 58 442
rect 68 444 86 446
rect 68 442 70 444
rect 72 442 82 444
rect 84 442 86 444
rect 68 440 86 442
rect 96 444 102 446
rect 96 442 98 444
rect 100 442 102 444
rect 96 440 102 442
rect 204 444 210 446
rect 204 442 206 444
rect 208 442 210 444
rect 204 440 210 442
rect 248 444 254 446
rect 248 442 250 444
rect 252 442 254 444
rect 248 440 254 442
rect 495 444 501 446
rect 495 442 497 444
rect 499 442 501 444
rect 495 440 501 442
rect 511 444 517 446
rect 511 442 513 444
rect 515 442 517 444
rect 511 440 517 442
rect 555 444 561 446
rect 555 442 557 444
rect 559 442 561 444
rect 555 440 561 442
rect 667 444 673 446
rect 667 442 669 444
rect 671 442 673 444
rect 667 440 673 442
rect 68 432 74 434
rect 68 430 70 432
rect 72 430 74 432
rect 68 428 74 430
rect 117 432 123 434
rect 117 430 119 432
rect 121 430 123 432
rect 117 428 123 430
rect 198 432 204 434
rect 198 430 200 432
rect 202 430 204 432
rect 198 428 204 430
rect 216 432 234 434
rect 216 430 218 432
rect 220 430 230 432
rect 232 430 234 432
rect 216 428 234 430
rect 244 432 250 434
rect 244 430 246 432
rect 248 430 250 432
rect 244 428 250 430
rect 288 432 294 434
rect 288 430 290 432
rect 292 430 294 432
rect 288 428 294 430
rect 446 432 452 434
rect 446 430 448 432
rect 450 430 452 432
rect 446 428 452 430
rect 463 432 481 434
rect 463 430 465 432
rect 467 430 477 432
rect 479 430 481 432
rect 463 428 481 430
rect 519 432 525 434
rect 519 430 521 432
rect 523 430 525 432
rect 519 428 525 430
rect 539 432 545 434
rect 539 430 541 432
rect 543 430 545 432
rect 539 428 545 430
rect 623 432 629 434
rect 623 430 625 432
rect 627 430 629 432
rect 623 428 629 430
rect 76 300 82 302
rect 76 298 78 300
rect 80 298 82 300
rect 76 296 82 298
rect 160 300 166 302
rect 160 298 162 300
rect 164 298 166 300
rect 160 296 166 298
rect 180 300 186 302
rect 180 298 182 300
rect 184 298 186 300
rect 180 296 186 298
rect 224 300 242 302
rect 224 298 226 300
rect 228 298 238 300
rect 240 298 242 300
rect 224 296 242 298
rect 253 300 259 302
rect 253 298 255 300
rect 257 298 259 300
rect 253 296 259 298
rect 411 300 417 302
rect 411 298 413 300
rect 415 298 417 300
rect 411 296 417 298
rect 455 300 461 302
rect 455 298 457 300
rect 459 298 461 300
rect 455 296 461 298
rect 471 300 489 302
rect 471 298 473 300
rect 475 298 485 300
rect 487 298 489 300
rect 471 296 489 298
rect 501 300 507 302
rect 501 298 503 300
rect 505 298 507 300
rect 501 296 507 298
rect 582 300 588 302
rect 582 298 584 300
rect 586 298 588 300
rect 582 296 588 298
rect 631 300 637 302
rect 631 298 633 300
rect 635 298 637 300
rect 631 296 637 298
rect 32 288 38 290
rect 32 286 34 288
rect 36 286 38 288
rect 32 284 38 286
rect 144 288 150 290
rect 144 286 146 288
rect 148 286 150 288
rect 144 284 150 286
rect 188 288 194 290
rect 188 286 190 288
rect 192 286 194 288
rect 188 284 194 286
rect 204 288 210 290
rect 204 286 206 288
rect 208 286 210 288
rect 204 284 210 286
rect 272 288 290 290
rect 272 286 274 288
rect 276 286 286 288
rect 288 286 290 288
rect 272 284 290 286
rect 451 288 457 290
rect 451 286 453 288
rect 455 286 457 288
rect 451 284 457 286
rect 495 288 501 290
rect 495 286 497 288
rect 499 286 501 288
rect 495 284 501 286
rect 603 288 609 290
rect 603 286 605 288
rect 607 286 609 288
rect 603 284 609 286
rect 619 288 637 290
rect 619 286 621 288
rect 623 286 633 288
rect 635 286 637 288
rect 619 284 637 286
rect 647 288 653 290
rect 647 286 649 288
rect 651 286 653 288
rect 647 284 653 286
rect 68 156 74 167
rect 68 154 70 156
rect 72 154 74 156
rect 68 152 74 154
rect 82 156 100 158
rect 82 154 84 156
rect 86 154 96 156
rect 98 154 100 156
rect 82 152 100 154
rect 112 156 118 158
rect 112 154 114 156
rect 116 154 118 156
rect 112 152 118 154
rect 192 156 198 167
rect 192 154 194 156
rect 196 154 198 156
rect 192 152 198 154
rect 447 156 453 158
rect 447 154 449 156
rect 451 154 453 156
rect 447 152 453 154
rect 555 156 561 173
rect 555 154 557 156
rect 559 154 561 156
rect 555 152 561 154
rect 667 156 673 158
rect 667 154 669 156
rect 671 154 673 156
rect 667 152 673 154
rect 32 144 38 146
rect 32 142 34 144
rect 36 142 38 144
rect 32 140 38 142
rect 166 144 172 146
rect 166 142 168 144
rect 170 142 172 144
rect 166 140 172 142
rect 186 144 204 146
rect 186 142 188 144
rect 190 142 200 144
rect 202 142 204 144
rect 186 140 204 142
rect 427 144 433 146
rect 427 142 429 144
rect 431 142 433 144
rect 427 125 433 142
rect 559 144 565 146
rect 559 142 561 144
rect 563 142 565 144
rect 559 140 565 142
rect 603 144 609 146
rect 603 142 605 144
rect 607 142 609 144
rect 603 140 609 142
rect 619 144 637 146
rect 619 142 621 144
rect 623 142 633 144
rect 635 142 637 144
rect 619 140 637 142
rect 68 12 74 23
rect 68 10 70 12
rect 72 10 74 12
rect 68 8 74 10
rect 80 12 98 14
rect 80 10 82 12
rect 84 10 94 12
rect 96 10 98 12
rect 80 8 98 10
rect 163 12 169 14
rect 163 10 165 12
rect 167 10 169 12
rect 163 8 169 10
rect 181 12 207 14
rect 181 10 183 12
rect 185 10 203 12
rect 205 10 207 12
rect 181 8 207 10
rect 377 12 395 14
rect 377 10 379 12
rect 381 10 391 12
rect 393 10 395 12
rect 377 8 395 10
rect 519 12 525 14
rect 519 10 521 12
rect 523 10 525 12
rect 519 8 525 10
rect 563 12 569 14
rect 563 10 565 12
rect 567 10 569 12
rect 563 8 569 10
rect 579 12 585 14
rect 579 10 581 12
rect 583 10 585 12
rect 579 8 585 10
rect 667 12 673 14
rect 667 10 669 12
rect 671 10 673 12
rect 667 8 673 10
<< ntie >>
rect 65 660 71 662
rect 65 658 67 660
rect 69 658 71 660
rect 136 660 142 662
rect 65 656 71 658
rect 136 658 138 660
rect 140 658 142 660
rect 213 660 219 662
rect 136 656 142 658
rect 213 658 215 660
rect 217 658 219 660
rect 213 656 219 658
rect 310 660 328 662
rect 517 660 523 662
rect 310 658 312 660
rect 314 658 324 660
rect 326 658 328 660
rect 310 656 328 658
rect 517 658 519 660
rect 521 658 523 660
rect 569 660 575 662
rect 517 656 523 658
rect 569 658 571 660
rect 573 658 575 660
rect 607 660 625 662
rect 569 656 575 658
rect 607 658 609 660
rect 611 658 621 660
rect 623 658 625 660
rect 607 656 625 658
rect 68 648 86 650
rect 68 646 70 648
rect 72 646 82 648
rect 84 646 86 648
rect 68 644 86 646
rect 96 648 102 650
rect 96 646 98 648
rect 100 646 102 648
rect 96 644 102 646
rect 184 648 190 650
rect 184 646 186 648
rect 188 646 190 648
rect 184 644 190 646
rect 250 648 278 650
rect 250 646 252 648
rect 254 646 274 648
rect 276 646 278 648
rect 250 644 278 646
rect 501 648 519 650
rect 501 646 503 648
rect 505 646 515 648
rect 517 646 519 648
rect 501 644 519 646
rect 533 648 539 650
rect 533 646 535 648
rect 537 646 539 648
rect 634 648 640 650
rect 533 644 539 646
rect 634 646 636 648
rect 638 646 640 648
rect 634 644 640 646
rect 65 516 71 518
rect 65 514 67 516
rect 69 514 71 516
rect 208 516 214 518
rect 65 512 71 514
rect 208 514 210 516
rect 212 514 214 516
rect 208 512 214 514
rect 443 516 461 518
rect 443 514 445 516
rect 447 514 457 516
rect 459 514 461 516
rect 587 516 593 518
rect 443 512 461 514
rect 587 514 589 516
rect 591 514 593 516
rect 587 512 593 514
rect 605 516 623 518
rect 605 514 607 516
rect 609 514 619 516
rect 621 514 623 516
rect 605 512 623 514
rect 68 504 86 506
rect 68 502 70 504
rect 72 502 82 504
rect 84 502 86 504
rect 68 500 86 502
rect 96 504 102 506
rect 96 502 98 504
rect 100 502 102 504
rect 171 504 177 506
rect 96 500 102 502
rect 171 502 173 504
rect 175 502 177 504
rect 248 504 254 506
rect 171 500 177 502
rect 248 502 250 504
rect 252 502 254 504
rect 462 504 468 506
rect 248 500 254 502
rect 462 502 464 504
rect 466 502 468 504
rect 511 504 517 506
rect 462 500 468 502
rect 511 502 513 504
rect 515 502 517 504
rect 511 500 517 502
rect 555 504 569 506
rect 555 502 557 504
rect 559 502 565 504
rect 567 502 569 504
rect 634 504 640 506
rect 555 500 569 502
rect 634 502 636 504
rect 638 502 640 504
rect 634 500 640 502
rect 33 372 47 374
rect 33 370 35 372
rect 37 370 43 372
rect 45 370 47 372
rect 33 368 47 370
rect 68 372 74 374
rect 68 370 70 372
rect 72 370 74 372
rect 68 368 74 370
rect 117 372 123 374
rect 117 370 119 372
rect 121 370 123 372
rect 117 368 123 370
rect 198 372 204 374
rect 198 370 200 372
rect 202 370 204 372
rect 198 368 204 370
rect 216 372 234 374
rect 216 370 218 372
rect 220 370 230 372
rect 232 370 234 372
rect 216 368 234 370
rect 244 372 250 374
rect 244 370 246 372
rect 248 370 250 372
rect 244 368 250 370
rect 332 372 338 374
rect 332 370 334 372
rect 336 370 338 372
rect 332 368 338 370
rect 446 372 452 374
rect 446 370 448 372
rect 450 370 452 372
rect 446 368 452 370
rect 463 372 481 374
rect 463 370 465 372
rect 467 370 477 372
rect 479 370 481 372
rect 463 368 481 370
rect 519 372 525 374
rect 519 370 521 372
rect 523 370 525 372
rect 519 368 525 370
rect 539 372 545 374
rect 539 370 541 372
rect 543 370 545 372
rect 539 368 545 370
rect 579 372 585 374
rect 579 370 581 372
rect 583 370 585 372
rect 579 368 585 370
rect 120 360 126 362
rect 120 358 122 360
rect 124 358 126 360
rect 120 356 126 358
rect 160 360 166 362
rect 160 358 162 360
rect 164 358 166 360
rect 160 356 166 358
rect 180 360 186 362
rect 180 358 182 360
rect 184 358 186 360
rect 180 356 186 358
rect 224 360 242 362
rect 224 358 226 360
rect 228 358 238 360
rect 240 358 242 360
rect 224 356 242 358
rect 253 360 259 362
rect 253 358 255 360
rect 257 358 259 360
rect 253 356 259 358
rect 367 360 373 362
rect 367 358 369 360
rect 371 358 373 360
rect 367 356 373 358
rect 455 360 461 362
rect 455 358 457 360
rect 459 358 461 360
rect 455 356 461 358
rect 471 360 489 362
rect 471 358 473 360
rect 475 358 485 360
rect 487 358 489 360
rect 471 356 489 358
rect 501 360 507 362
rect 501 358 503 360
rect 505 358 507 360
rect 501 356 507 358
rect 582 360 588 362
rect 582 358 584 360
rect 586 358 588 360
rect 582 356 588 358
rect 631 360 637 362
rect 631 358 633 360
rect 635 358 637 360
rect 631 356 637 358
rect 658 360 672 362
rect 658 358 660 360
rect 662 358 668 360
rect 670 358 672 360
rect 658 356 672 358
rect 65 228 71 230
rect 65 226 67 228
rect 69 226 71 228
rect 136 228 150 230
rect 65 224 71 226
rect 136 226 138 228
rect 140 226 146 228
rect 148 226 150 228
rect 136 224 150 226
rect 188 228 194 230
rect 188 226 190 228
rect 192 226 194 228
rect 237 228 243 230
rect 188 224 194 226
rect 237 226 239 228
rect 241 226 243 228
rect 272 228 290 230
rect 237 224 243 226
rect 272 226 274 228
rect 276 226 286 228
rect 288 226 290 228
rect 272 224 290 226
rect 451 228 457 230
rect 451 226 453 228
rect 455 226 457 228
rect 528 228 534 230
rect 451 224 457 226
rect 528 226 530 228
rect 532 226 534 228
rect 603 228 609 230
rect 528 224 534 226
rect 603 226 605 228
rect 607 226 609 228
rect 603 224 609 226
rect 619 228 637 230
rect 619 226 621 228
rect 623 226 633 228
rect 635 226 637 228
rect 619 224 637 226
rect 82 216 100 218
rect 82 214 84 216
rect 86 214 96 216
rect 98 214 100 216
rect 82 212 100 214
rect 112 216 118 218
rect 112 214 114 216
rect 116 214 118 216
rect 112 212 118 214
rect 491 216 497 218
rect 491 214 493 216
rect 495 214 497 216
rect 634 216 640 218
rect 491 212 497 214
rect 634 214 636 216
rect 638 214 640 216
rect 634 212 640 214
rect 65 84 71 86
rect 65 82 67 84
rect 69 82 71 84
rect 166 84 172 86
rect 65 80 71 82
rect 166 82 168 84
rect 170 82 172 84
rect 166 80 172 82
rect 186 84 204 86
rect 186 82 188 84
rect 190 82 200 84
rect 202 82 204 84
rect 186 80 204 82
rect 427 84 455 86
rect 427 82 429 84
rect 431 82 451 84
rect 453 82 455 84
rect 427 80 455 82
rect 515 84 521 86
rect 515 82 517 84
rect 519 82 521 84
rect 515 80 521 82
rect 603 84 609 86
rect 603 82 605 84
rect 607 82 609 84
rect 603 80 609 82
rect 619 84 637 86
rect 619 82 621 84
rect 623 82 633 84
rect 635 82 637 84
rect 619 80 637 82
rect 80 72 98 74
rect 80 70 82 72
rect 84 70 94 72
rect 96 70 98 72
rect 130 72 136 74
rect 80 68 98 70
rect 130 70 132 72
rect 134 70 136 72
rect 182 72 188 74
rect 130 68 136 70
rect 182 70 184 72
rect 186 70 188 72
rect 377 72 395 74
rect 377 70 379 72
rect 381 70 391 72
rect 393 70 395 72
rect 182 68 188 70
rect 377 68 395 70
rect 486 72 492 74
rect 486 70 488 72
rect 490 70 492 72
rect 563 72 569 74
rect 486 68 492 70
rect 563 70 565 72
rect 567 70 569 72
rect 634 72 640 74
rect 563 68 569 70
rect 634 70 636 72
rect 638 70 640 72
rect 634 68 640 70
<< nmos >>
rect 38 699 40 708
rect 54 704 56 713
rect 64 704 66 713
rect 74 704 76 716
rect 81 704 83 716
rect 107 705 109 713
rect 118 702 120 710
rect 142 701 144 710
rect 155 701 157 712
rect 162 701 164 712
rect 186 699 188 708
rect 202 704 204 713
rect 212 704 214 713
rect 222 704 224 716
rect 229 704 231 716
rect 262 699 264 719
rect 269 699 271 719
rect 276 699 278 719
rect 283 699 285 719
rect 316 699 318 708
rect 505 699 507 709
rect 515 699 517 709
rect 542 699 544 708
rect 558 704 560 713
rect 568 704 570 713
rect 578 704 580 716
rect 585 704 587 716
rect 613 699 615 708
rect 653 704 655 719
rect 663 704 665 719
rect 41 587 43 607
rect 48 587 50 607
rect 74 598 76 607
rect 102 596 104 605
rect 115 594 117 605
rect 122 594 124 605
rect 146 597 148 606
rect 159 593 161 606
rect 166 593 168 606
rect 173 593 175 606
rect 214 593 216 599
rect 224 593 226 599
rect 236 593 238 599
rect 246 593 248 599
rect 511 598 513 607
rect 539 596 541 605
rect 552 594 554 605
rect 559 594 561 605
rect 587 587 589 607
rect 594 587 596 607
rect 622 590 624 602
rect 629 590 631 602
rect 639 593 641 602
rect 649 593 651 602
rect 665 598 667 607
rect 38 555 40 564
rect 54 560 56 569
rect 64 560 66 569
rect 74 560 76 572
rect 81 560 83 572
rect 109 555 111 575
rect 116 555 118 575
rect 168 563 170 573
rect 178 563 180 573
rect 190 563 192 573
rect 223 556 225 569
rect 230 556 232 569
rect 237 556 239 569
rect 250 556 252 565
rect 449 555 451 564
rect 529 560 531 575
rect 539 560 541 575
rect 565 557 567 568
rect 572 557 574 568
rect 585 557 587 566
rect 611 555 613 564
rect 653 560 655 575
rect 663 560 665 575
rect 39 449 41 457
rect 50 452 52 460
rect 74 454 76 463
rect 102 452 104 461
rect 115 450 117 461
rect 122 450 124 461
rect 159 446 161 458
rect 166 446 168 458
rect 176 449 178 458
rect 186 449 188 458
rect 202 454 204 463
rect 226 450 228 461
rect 233 450 235 461
rect 246 452 248 461
rect 450 446 452 458
rect 457 446 459 458
rect 467 449 469 458
rect 477 449 479 458
rect 493 454 495 463
rect 517 452 519 461
rect 530 450 532 461
rect 537 450 539 461
rect 561 452 563 463
rect 572 444 574 463
rect 582 448 584 463
rect 592 448 594 463
rect 622 446 624 458
rect 629 446 631 458
rect 639 449 641 458
rect 649 449 651 458
rect 665 454 667 463
rect 44 418 46 430
rect 51 418 53 430
rect 74 413 76 422
rect 87 413 89 424
rect 94 413 96 424
rect 123 413 125 422
rect 136 413 138 424
rect 143 413 145 424
rect 176 413 178 424
rect 183 413 185 424
rect 196 413 198 422
rect 222 411 224 420
rect 250 413 252 422
rect 263 413 265 424
rect 270 413 272 424
rect 294 412 296 421
rect 307 412 309 425
rect 314 412 316 425
rect 321 412 323 425
rect 424 413 426 424
rect 431 413 433 424
rect 444 413 446 422
rect 469 411 471 420
rect 497 413 499 424
rect 504 413 506 424
rect 517 413 519 422
rect 545 413 547 422
rect 558 413 560 424
rect 565 413 567 424
rect 594 412 596 425
rect 601 412 603 425
rect 608 412 610 425
rect 621 412 623 421
rect 648 411 650 431
rect 655 411 657 431
rect 662 411 664 431
rect 41 299 43 319
rect 48 299 50 319
rect 55 299 57 319
rect 82 309 84 318
rect 95 305 97 318
rect 102 305 104 318
rect 109 305 111 318
rect 138 306 140 317
rect 145 306 147 317
rect 158 308 160 317
rect 186 308 188 317
rect 199 306 201 317
rect 206 306 208 317
rect 234 310 236 319
rect 259 308 261 317
rect 272 306 274 317
rect 279 306 281 317
rect 382 305 384 318
rect 389 305 391 318
rect 396 305 398 318
rect 409 309 411 318
rect 433 306 435 317
rect 440 306 442 317
rect 453 308 455 317
rect 481 310 483 319
rect 507 308 509 317
rect 520 306 522 317
rect 527 306 529 317
rect 560 306 562 317
rect 567 306 569 317
rect 580 308 582 317
rect 609 306 611 317
rect 616 306 618 317
rect 629 308 631 317
rect 652 300 654 312
rect 659 300 661 312
rect 38 267 40 276
rect 54 272 56 281
rect 64 272 66 281
rect 74 272 76 284
rect 81 272 83 284
rect 111 267 113 282
rect 121 267 123 282
rect 131 267 133 286
rect 142 267 144 278
rect 166 269 168 280
rect 173 269 175 280
rect 186 269 188 278
rect 210 267 212 276
rect 226 272 228 281
rect 236 272 238 281
rect 246 272 248 284
rect 253 272 255 284
rect 278 267 280 276
rect 457 269 459 278
rect 470 269 472 280
rect 477 269 479 280
rect 501 267 503 276
rect 517 272 519 281
rect 527 272 529 281
rect 537 272 539 284
rect 544 272 546 284
rect 581 269 583 280
rect 588 269 590 280
rect 601 269 603 278
rect 629 267 631 276
rect 653 270 655 278
rect 664 273 666 281
rect 40 155 42 170
rect 50 155 52 170
rect 92 166 94 175
rect 118 164 120 173
rect 131 162 133 173
rect 138 162 140 173
rect 164 155 166 170
rect 174 155 176 170
rect 453 165 455 174
rect 466 161 468 174
rect 473 161 475 174
rect 480 161 482 174
rect 513 157 515 167
rect 525 157 527 167
rect 535 157 537 167
rect 587 155 589 175
rect 594 155 596 175
rect 622 158 624 170
rect 629 158 631 170
rect 639 161 641 170
rect 649 161 651 170
rect 665 166 667 175
rect 38 123 40 132
rect 54 128 56 137
rect 64 128 66 137
rect 74 128 76 140
rect 81 128 83 140
rect 109 123 111 143
rect 116 123 118 143
rect 144 125 146 136
rect 151 125 153 136
rect 164 125 166 134
rect 192 123 194 132
rect 457 131 459 137
rect 467 131 469 137
rect 479 131 481 137
rect 489 131 491 137
rect 530 124 532 137
rect 537 124 539 137
rect 544 124 546 137
rect 557 124 559 133
rect 581 125 583 136
rect 588 125 590 136
rect 601 125 603 134
rect 629 123 631 132
rect 655 123 657 143
rect 662 123 664 143
rect 40 11 42 26
rect 50 11 52 26
rect 90 22 92 31
rect 118 14 120 26
rect 125 14 127 26
rect 135 17 137 26
rect 145 17 147 26
rect 161 22 163 31
rect 188 21 190 31
rect 198 21 200 31
rect 387 22 389 31
rect 420 11 422 31
rect 427 11 429 31
rect 434 11 436 31
rect 441 11 443 31
rect 474 14 476 26
rect 481 14 483 26
rect 491 17 493 26
rect 501 17 503 26
rect 517 22 519 31
rect 541 18 543 29
rect 548 18 550 29
rect 561 20 563 29
rect 585 20 587 28
rect 596 17 598 25
rect 622 14 624 26
rect 629 14 631 26
rect 639 17 641 26
rect 649 17 651 26
rect 665 22 667 31
<< pmos >>
rect 46 659 48 686
rect 62 668 64 686
rect 72 668 74 686
rect 82 659 84 686
rect 109 659 111 687
rect 116 659 118 687
rect 142 668 144 686
rect 152 666 154 679
rect 162 666 164 679
rect 194 659 196 686
rect 210 668 212 686
rect 220 668 222 686
rect 230 659 232 686
rect 256 663 258 680
rect 266 663 268 680
rect 276 663 278 680
rect 286 663 288 680
rect 316 669 318 687
rect 505 660 507 684
rect 515 668 517 684
rect 550 659 552 686
rect 566 668 568 686
rect 576 668 578 686
rect 586 659 588 686
rect 613 669 615 687
rect 641 659 643 686
rect 648 659 650 686
rect 658 659 660 686
rect 665 659 667 686
rect 38 623 40 647
rect 48 623 50 647
rect 74 619 76 637
rect 102 620 104 638
rect 112 627 114 640
rect 122 627 124 640
rect 146 621 148 639
rect 156 626 158 639
rect 166 626 168 639
rect 178 625 180 638
rect 218 620 220 645
rect 225 620 227 645
rect 232 620 234 645
rect 239 620 241 645
rect 249 620 251 638
rect 256 620 258 638
rect 263 620 265 638
rect 270 620 272 638
rect 511 619 513 637
rect 539 620 541 638
rect 549 627 551 640
rect 559 627 561 640
rect 587 623 589 647
rect 597 623 599 647
rect 621 620 623 647
rect 631 620 633 638
rect 641 620 643 638
rect 657 620 659 647
rect 46 515 48 542
rect 62 524 64 542
rect 72 524 74 542
rect 82 515 84 542
rect 106 515 108 539
rect 116 515 118 539
rect 150 515 152 543
rect 157 515 159 543
rect 164 515 166 543
rect 174 515 176 543
rect 181 515 183 543
rect 188 515 190 543
rect 218 524 220 537
rect 230 523 232 536
rect 240 523 242 536
rect 250 523 252 541
rect 449 525 451 543
rect 517 515 519 542
rect 524 515 526 542
rect 534 515 536 542
rect 541 515 543 542
rect 565 522 567 535
rect 575 522 577 535
rect 585 524 587 542
rect 611 525 613 543
rect 641 515 643 542
rect 648 515 650 542
rect 658 515 660 542
rect 665 515 667 542
rect 41 475 43 503
rect 48 475 50 503
rect 74 475 76 493
rect 102 476 104 494
rect 112 483 114 496
rect 122 483 124 496
rect 158 476 160 503
rect 168 476 170 494
rect 178 476 180 494
rect 194 476 196 503
rect 226 483 228 496
rect 236 483 238 496
rect 246 476 248 494
rect 449 476 451 503
rect 459 476 461 494
rect 469 476 471 494
rect 485 476 487 503
rect 517 476 519 494
rect 527 483 529 496
rect 537 483 539 496
rect 562 476 564 494
rect 572 476 574 494
rect 582 476 584 494
rect 592 476 594 494
rect 621 476 623 503
rect 631 476 633 494
rect 641 476 643 494
rect 657 476 659 503
rect 40 380 42 394
rect 50 380 52 394
rect 74 380 76 398
rect 84 378 86 391
rect 94 378 96 391
rect 123 380 125 398
rect 133 378 135 391
rect 143 378 145 391
rect 176 378 178 391
rect 186 378 188 391
rect 196 380 198 398
rect 222 381 224 399
rect 250 380 252 398
rect 260 378 262 391
rect 270 378 272 391
rect 294 379 296 397
rect 304 379 306 392
rect 314 379 316 392
rect 326 380 328 393
rect 424 378 426 391
rect 434 378 436 391
rect 444 380 446 398
rect 469 381 471 399
rect 497 378 499 391
rect 507 378 509 391
rect 517 380 519 398
rect 545 380 547 398
rect 555 378 557 391
rect 565 378 567 391
rect 589 380 591 393
rect 601 379 603 392
rect 611 379 613 392
rect 621 379 623 397
rect 645 371 647 391
rect 655 371 657 391
rect 665 371 667 391
rect 38 339 40 359
rect 48 339 50 359
rect 58 339 60 359
rect 82 333 84 351
rect 92 338 94 351
rect 102 338 104 351
rect 114 337 116 350
rect 138 339 140 352
rect 148 339 150 352
rect 158 332 160 350
rect 186 332 188 350
rect 196 339 198 352
rect 206 339 208 352
rect 234 331 236 349
rect 259 332 261 350
rect 269 339 271 352
rect 279 339 281 352
rect 377 337 379 350
rect 389 338 391 351
rect 399 338 401 351
rect 409 333 411 351
rect 433 339 435 352
rect 443 339 445 352
rect 453 332 455 350
rect 481 331 483 349
rect 507 332 509 350
rect 517 339 519 352
rect 527 339 529 352
rect 560 339 562 352
rect 570 339 572 352
rect 580 332 582 350
rect 609 339 611 352
rect 619 339 621 352
rect 629 332 631 350
rect 653 336 655 350
rect 663 336 665 350
rect 46 227 48 254
rect 62 236 64 254
rect 72 236 74 254
rect 82 227 84 254
rect 111 236 113 254
rect 121 236 123 254
rect 131 236 133 254
rect 141 236 143 254
rect 166 234 168 247
rect 176 234 178 247
rect 186 236 188 254
rect 218 227 220 254
rect 234 236 236 254
rect 244 236 246 254
rect 254 227 256 254
rect 278 237 280 255
rect 457 236 459 254
rect 467 234 469 247
rect 477 234 479 247
rect 509 227 511 254
rect 525 236 527 254
rect 535 236 537 254
rect 545 227 547 254
rect 581 234 583 247
rect 591 234 593 247
rect 601 236 603 254
rect 629 237 631 255
rect 655 227 657 255
rect 662 227 664 255
rect 38 188 40 215
rect 45 188 47 215
rect 55 188 57 215
rect 62 188 64 215
rect 92 187 94 205
rect 118 188 120 206
rect 128 195 130 208
rect 138 195 140 208
rect 162 188 164 215
rect 169 188 171 215
rect 179 188 181 215
rect 186 188 188 215
rect 453 189 455 207
rect 463 194 465 207
rect 473 194 475 207
rect 485 193 487 206
rect 515 187 517 215
rect 522 187 524 215
rect 529 187 531 215
rect 539 187 541 215
rect 546 187 548 215
rect 553 187 555 215
rect 587 191 589 215
rect 597 191 599 215
rect 621 188 623 215
rect 631 188 633 206
rect 641 188 643 206
rect 657 188 659 215
rect 46 83 48 110
rect 62 92 64 110
rect 72 92 74 110
rect 82 83 84 110
rect 106 83 108 107
rect 116 83 118 107
rect 144 90 146 103
rect 154 90 156 103
rect 164 92 166 110
rect 192 93 194 111
rect 433 92 435 110
rect 440 92 442 110
rect 447 92 449 110
rect 454 92 456 110
rect 464 85 466 110
rect 471 85 473 110
rect 478 85 480 110
rect 485 85 487 110
rect 525 92 527 105
rect 537 91 539 104
rect 547 91 549 104
rect 557 91 559 109
rect 581 90 583 103
rect 591 90 593 103
rect 601 92 603 110
rect 629 93 631 111
rect 655 83 657 107
rect 665 83 667 107
rect 38 44 40 71
rect 45 44 47 71
rect 55 44 57 71
rect 62 44 64 71
rect 90 43 92 61
rect 117 44 119 71
rect 127 44 129 62
rect 137 44 139 62
rect 153 44 155 71
rect 188 46 190 62
rect 198 46 200 70
rect 387 43 389 61
rect 417 50 419 67
rect 427 50 429 67
rect 437 50 439 67
rect 447 50 449 67
rect 473 44 475 71
rect 483 44 485 62
rect 493 44 495 62
rect 509 44 511 71
rect 541 51 543 64
rect 551 51 553 64
rect 561 44 563 62
rect 587 43 589 71
rect 594 43 596 71
rect 621 44 623 71
rect 631 44 633 62
rect 641 44 643 62
rect 657 44 659 71
<< polyct0 >>
rect 70 692 72 694
rect 80 691 82 693
rect 144 692 146 694
rect 218 692 220 694
rect 228 691 230 693
rect 574 692 576 694
rect 278 685 280 687
rect 584 691 586 693
rect 104 612 106 614
rect 148 612 150 614
rect 541 612 543 614
rect 623 613 625 615
rect 633 612 635 614
rect 70 548 72 550
rect 80 547 82 549
rect 248 548 250 550
rect 583 548 585 550
rect 104 468 106 470
rect 160 469 162 471
rect 170 468 172 470
rect 244 468 246 470
rect 451 469 453 471
rect 461 468 463 470
rect 519 468 521 470
rect 623 469 625 471
rect 633 468 635 470
rect 76 404 78 406
rect 125 404 127 406
rect 194 404 196 406
rect 252 404 254 406
rect 296 404 298 406
rect 442 404 444 406
rect 515 404 517 406
rect 547 404 549 406
rect 619 404 621 406
rect 84 324 86 326
rect 156 324 158 326
rect 188 324 190 326
rect 261 324 263 326
rect 407 324 409 326
rect 451 324 453 326
rect 509 324 511 326
rect 578 324 580 326
rect 627 324 629 326
rect 70 260 72 262
rect 80 259 82 261
rect 184 260 186 262
rect 242 260 244 262
rect 252 259 254 261
rect 459 260 461 262
rect 533 260 535 262
rect 543 259 545 261
rect 599 260 601 262
rect 120 180 122 182
rect 455 180 457 182
rect 623 181 625 183
rect 633 180 635 182
rect 70 116 72 118
rect 80 115 82 117
rect 162 116 164 118
rect 555 116 557 118
rect 599 116 601 118
rect 119 37 121 39
rect 425 43 427 45
rect 129 36 131 38
rect 475 37 477 39
rect 485 36 487 38
rect 559 36 561 38
rect 623 37 625 39
rect 633 36 635 38
<< polyct1 >>
rect 49 697 51 699
rect 108 692 110 694
rect 118 695 120 697
rect 154 692 156 694
rect 33 684 35 686
rect 197 697 199 699
rect 164 684 166 686
rect 258 692 260 694
rect 181 684 183 686
rect 290 692 292 694
rect 318 692 320 694
rect 521 691 523 693
rect 553 697 555 699
rect 639 700 641 702
rect 268 685 270 687
rect 615 692 617 694
rect 537 684 539 686
rect 661 697 663 699
rect 650 692 652 694
rect 55 616 57 618
rect 40 612 42 614
rect 124 620 126 622
rect 76 612 78 614
rect 114 612 116 614
rect 168 619 170 621
rect 158 612 160 614
rect 180 612 182 614
rect 209 613 211 615
rect 224 606 226 608
rect 235 604 237 606
rect 274 613 276 615
rect 509 612 511 614
rect 254 604 256 606
rect 264 607 266 609
rect 561 620 563 622
rect 551 612 553 614
rect 264 596 266 598
rect 580 616 582 618
rect 670 620 672 622
rect 595 612 597 614
rect 654 607 656 609
rect 49 553 51 555
rect 108 548 110 550
rect 155 554 157 556
rect 145 548 147 550
rect 33 540 35 542
rect 123 544 125 546
rect 166 556 168 558
rect 178 556 180 558
rect 188 556 190 558
rect 216 548 218 550
rect 515 556 517 558
rect 238 548 240 550
rect 228 541 230 543
rect 451 548 453 550
rect 537 553 539 555
rect 526 548 528 550
rect 639 556 641 558
rect 573 548 575 550
rect 563 540 565 542
rect 613 548 615 550
rect 661 553 663 555
rect 650 548 652 550
rect 40 468 42 470
rect 124 476 126 478
rect 207 476 209 478
rect 50 465 52 467
rect 76 468 78 470
rect 114 468 116 470
rect 224 476 226 478
rect 191 463 193 465
rect 498 476 500 478
rect 234 468 236 470
rect 539 476 541 478
rect 670 476 672 478
rect 482 463 484 465
rect 529 468 531 470
rect 563 468 565 470
rect 595 468 597 470
rect 654 463 656 465
rect 38 411 40 413
rect 49 404 51 406
rect 86 404 88 406
rect 135 404 137 406
rect 96 396 98 398
rect 184 404 186 406
rect 145 396 147 398
rect 174 396 176 398
rect 224 404 226 406
rect 262 404 264 406
rect 306 404 308 406
rect 272 396 274 398
rect 328 404 330 406
rect 316 397 318 399
rect 432 404 434 406
rect 422 396 424 398
rect 471 404 473 406
rect 505 404 507 406
rect 495 396 497 398
rect 557 404 559 406
rect 587 404 589 406
rect 567 396 569 398
rect 609 404 611 406
rect 643 404 645 406
rect 599 397 601 399
rect 663 404 665 406
rect 653 396 655 398
rect 50 332 52 334
rect 40 324 42 326
rect 104 331 106 333
rect 60 324 62 326
rect 94 324 96 326
rect 136 332 138 334
rect 116 324 118 326
rect 146 324 148 326
rect 208 332 210 334
rect 198 324 200 326
rect 232 324 234 326
rect 281 332 283 334
rect 271 324 273 326
rect 387 331 389 333
rect 375 324 377 326
rect 431 332 433 334
rect 397 324 399 326
rect 441 324 443 326
rect 479 324 481 326
rect 529 332 531 334
rect 558 332 560 334
rect 519 324 521 326
rect 607 332 609 334
rect 568 324 570 326
rect 617 324 619 326
rect 654 324 656 326
rect 665 317 667 319
rect 49 265 51 267
rect 108 260 110 262
rect 140 260 142 262
rect 174 260 176 262
rect 221 265 223 267
rect 33 252 35 254
rect 164 252 166 254
rect 280 260 282 262
rect 469 260 471 262
rect 205 252 207 254
rect 512 265 514 267
rect 479 252 481 254
rect 589 260 591 262
rect 627 260 629 262
rect 653 263 655 265
rect 496 252 498 254
rect 579 252 581 254
rect 663 260 665 262
rect 53 180 55 182
rect 42 175 44 177
rect 90 180 92 182
rect 140 188 142 190
rect 130 180 132 182
rect 64 172 66 174
rect 177 180 179 182
rect 166 175 168 177
rect 475 187 477 189
rect 465 180 467 182
rect 487 180 489 182
rect 188 172 190 174
rect 515 172 517 174
rect 525 172 527 174
rect 537 172 539 174
rect 580 184 582 186
rect 670 188 672 190
rect 558 180 560 182
rect 548 174 550 176
rect 595 180 597 182
rect 654 175 656 177
rect 49 121 51 123
rect 108 116 110 118
rect 33 108 35 110
rect 123 112 125 114
rect 439 132 441 134
rect 152 116 154 118
rect 142 108 144 110
rect 439 121 441 123
rect 449 124 451 126
rect 194 116 196 118
rect 429 115 431 117
rect 468 124 470 126
rect 479 122 481 124
rect 494 115 496 117
rect 523 116 525 118
rect 545 116 547 118
rect 535 109 537 111
rect 589 116 591 118
rect 627 116 629 118
rect 579 108 581 110
rect 663 116 665 118
rect 648 112 650 114
rect 53 36 55 38
rect 42 31 44 33
rect 166 44 168 46
rect 88 36 90 38
rect 435 43 437 45
rect 64 28 66 30
rect 150 31 152 33
rect 182 37 184 39
rect 385 36 387 38
rect 413 36 415 38
rect 522 44 524 46
rect 445 36 447 38
rect 539 44 541 46
rect 506 31 508 33
rect 670 44 672 46
rect 549 36 551 38
rect 585 33 587 35
rect 595 36 597 38
rect 654 31 656 33
<< ndifct0 >>
rect 47 709 49 711
rect 33 701 35 703
rect 59 706 61 708
rect 123 706 125 708
rect 167 708 169 710
rect 195 709 197 711
rect 181 701 183 703
rect 207 706 209 708
rect 499 708 501 710
rect 325 704 327 706
rect 551 709 553 711
rect 521 705 523 707
rect 537 701 539 703
rect 563 706 565 708
rect 648 715 650 717
rect 648 708 650 710
rect 622 704 624 706
rect 668 715 670 717
rect 83 600 85 602
rect 55 596 57 598
rect 127 596 129 598
rect 55 589 57 591
rect 178 595 180 597
rect 209 595 211 597
rect 251 595 253 597
rect 502 600 504 602
rect 564 596 566 598
rect 580 596 582 598
rect 580 589 582 591
rect 644 598 646 600
rect 670 603 672 605
rect 656 595 658 597
rect 47 565 49 567
rect 33 557 35 559
rect 59 562 61 564
rect 123 571 125 573
rect 123 564 125 566
rect 218 565 220 567
rect 524 571 526 573
rect 524 564 526 566
rect 458 560 460 562
rect 544 571 546 573
rect 560 564 562 566
rect 648 571 650 573
rect 648 564 650 566
rect 620 560 622 562
rect 668 571 670 573
rect 55 454 57 456
rect 83 456 85 458
rect 127 452 129 454
rect 181 454 183 456
rect 207 459 209 461
rect 193 451 195 453
rect 221 452 223 454
rect 472 454 474 456
rect 498 459 500 461
rect 484 451 486 453
rect 556 459 558 461
rect 542 452 544 454
rect 567 450 569 452
rect 577 458 579 460
rect 577 451 579 453
rect 597 451 599 453
rect 644 454 646 456
rect 670 459 672 461
rect 656 451 658 453
rect 34 426 36 428
rect 99 420 101 422
rect 148 420 150 422
rect 171 420 173 422
rect 231 416 233 418
rect 275 420 277 422
rect 326 421 328 423
rect 419 420 421 422
rect 492 420 494 422
rect 478 416 480 418
rect 642 428 644 429
rect 570 420 572 422
rect 589 421 591 423
rect 114 307 116 309
rect 133 308 135 310
rect 61 301 63 302
rect 225 312 227 314
rect 211 308 213 310
rect 284 308 286 310
rect 377 307 379 309
rect 428 308 430 310
rect 472 312 474 314
rect 532 308 534 310
rect 555 308 557 310
rect 604 308 606 310
rect 669 302 671 304
rect 47 277 49 279
rect 33 269 35 271
rect 59 274 61 276
rect 106 277 108 279
rect 126 277 128 279
rect 126 270 128 272
rect 136 278 138 280
rect 161 276 163 278
rect 147 269 149 271
rect 219 277 221 279
rect 205 269 207 271
rect 231 274 233 276
rect 287 272 289 274
rect 482 276 484 278
rect 510 277 512 279
rect 496 269 498 271
rect 522 274 524 276
rect 576 276 578 278
rect 620 272 622 274
rect 648 274 650 276
rect 35 157 37 159
rect 83 168 85 170
rect 55 164 57 166
rect 55 157 57 159
rect 143 164 145 166
rect 159 157 161 159
rect 179 164 181 166
rect 179 157 181 159
rect 485 163 487 165
rect 580 164 582 166
rect 580 157 582 159
rect 644 166 646 168
rect 670 171 672 173
rect 656 163 658 165
rect 47 133 49 135
rect 33 125 35 127
rect 59 130 61 132
rect 123 139 125 141
rect 123 132 125 134
rect 139 132 141 134
rect 201 128 203 130
rect 452 133 454 135
rect 494 133 496 135
rect 525 133 527 135
rect 648 139 650 141
rect 576 132 578 134
rect 648 132 650 134
rect 620 128 622 130
rect 35 13 37 15
rect 81 24 83 26
rect 55 20 57 22
rect 55 13 57 15
rect 140 22 142 24
rect 166 27 168 29
rect 182 23 184 25
rect 152 19 154 21
rect 378 24 380 26
rect 204 20 206 22
rect 496 22 498 24
rect 522 27 524 29
rect 508 19 510 21
rect 536 20 538 22
rect 580 22 582 24
rect 644 22 646 24
rect 670 27 672 29
rect 656 19 658 21
<< ndifct1 >>
rect 87 718 89 720
rect 69 708 71 710
rect 101 718 103 720
rect 148 718 150 720
rect 112 709 114 711
rect 235 718 237 720
rect 137 706 139 708
rect 217 708 219 710
rect 257 709 259 711
rect 289 718 291 720
rect 591 718 593 720
rect 311 701 313 703
rect 510 701 512 703
rect 573 708 575 710
rect 608 701 610 703
rect 658 708 660 710
rect 36 595 38 597
rect 69 603 71 605
rect 97 598 99 600
rect 141 602 143 604
rect 219 595 221 597
rect 241 595 243 597
rect 108 586 110 588
rect 516 603 518 605
rect 534 598 536 600
rect 152 586 154 588
rect 230 586 232 588
rect 545 586 547 588
rect 599 595 601 597
rect 634 596 636 598
rect 616 586 618 588
rect 87 574 89 576
rect 69 564 71 566
rect 104 565 106 567
rect 162 574 164 576
rect 184 574 186 576
rect 244 574 246 576
rect 173 565 175 567
rect 195 565 197 567
rect 255 558 257 560
rect 444 557 446 559
rect 534 564 536 566
rect 579 574 581 576
rect 590 562 592 564
rect 606 557 608 559
rect 658 564 660 566
rect 44 451 46 453
rect 69 459 71 461
rect 97 454 99 456
rect 33 442 35 444
rect 171 452 173 454
rect 251 454 253 456
rect 108 442 110 444
rect 153 442 155 444
rect 462 452 464 454
rect 512 454 514 456
rect 240 442 242 444
rect 444 442 446 444
rect 523 442 525 444
rect 587 459 589 461
rect 634 452 636 454
rect 616 442 618 444
rect 80 430 82 432
rect 129 430 131 432
rect 56 420 58 422
rect 69 418 71 420
rect 190 430 192 432
rect 256 430 258 432
rect 118 418 120 420
rect 300 430 302 432
rect 438 430 440 432
rect 201 418 203 420
rect 217 413 219 415
rect 245 418 247 420
rect 289 414 291 416
rect 511 430 513 432
rect 551 430 553 432
rect 615 430 617 432
rect 449 418 451 420
rect 464 413 466 415
rect 642 429 644 430
rect 522 418 524 420
rect 540 418 542 420
rect 626 414 628 416
rect 667 421 669 423
rect 36 307 38 309
rect 77 314 79 316
rect 163 310 165 312
rect 181 310 183 312
rect 61 300 63 301
rect 239 315 241 317
rect 254 310 256 312
rect 88 298 90 300
rect 152 298 154 300
rect 192 298 194 300
rect 414 314 416 316
rect 458 310 460 312
rect 486 315 488 317
rect 502 310 504 312
rect 265 298 267 300
rect 403 298 405 300
rect 585 310 587 312
rect 447 298 449 300
rect 513 298 515 300
rect 634 310 636 312
rect 647 308 649 310
rect 574 298 576 300
rect 623 298 625 300
rect 87 286 89 288
rect 69 276 71 278
rect 116 269 118 271
rect 180 286 182 288
rect 259 286 261 288
rect 463 286 465 288
rect 191 274 193 276
rect 241 276 243 278
rect 550 286 552 288
rect 595 286 597 288
rect 273 269 275 271
rect 452 274 454 276
rect 532 276 534 278
rect 670 286 672 288
rect 606 274 608 276
rect 634 269 636 271
rect 659 277 661 279
rect 45 164 47 166
rect 97 171 99 173
rect 113 166 115 168
rect 448 170 450 172
rect 124 154 126 156
rect 169 164 171 166
rect 508 163 510 165
rect 530 163 532 165
rect 459 154 461 156
rect 519 154 521 156
rect 541 154 543 156
rect 599 163 601 165
rect 634 164 636 166
rect 616 154 618 156
rect 87 142 89 144
rect 69 132 71 134
rect 104 133 106 135
rect 158 142 160 144
rect 473 142 475 144
rect 551 142 553 144
rect 169 130 171 132
rect 187 125 189 127
rect 595 142 597 144
rect 462 133 464 135
rect 484 133 486 135
rect 562 126 564 128
rect 606 130 608 132
rect 634 125 636 127
rect 667 133 669 135
rect 45 20 47 22
rect 95 27 97 29
rect 130 20 132 22
rect 193 27 195 29
rect 392 27 394 29
rect 112 10 114 12
rect 414 10 416 12
rect 446 19 448 21
rect 486 20 488 22
rect 566 22 568 24
rect 468 10 470 12
rect 591 19 593 21
rect 555 10 557 12
rect 602 10 604 12
rect 634 20 636 22
rect 616 10 618 12
<< ntiect1 >>
rect 67 658 69 660
rect 138 658 140 660
rect 215 658 217 660
rect 312 658 314 660
rect 324 658 326 660
rect 519 658 521 660
rect 571 658 573 660
rect 609 658 611 660
rect 621 658 623 660
rect 70 646 72 648
rect 82 646 84 648
rect 98 646 100 648
rect 186 646 188 648
rect 252 646 254 648
rect 274 646 276 648
rect 503 646 505 648
rect 515 646 517 648
rect 535 646 537 648
rect 636 646 638 648
rect 67 514 69 516
rect 210 514 212 516
rect 445 514 447 516
rect 457 514 459 516
rect 589 514 591 516
rect 607 514 609 516
rect 619 514 621 516
rect 70 502 72 504
rect 82 502 84 504
rect 98 502 100 504
rect 173 502 175 504
rect 250 502 252 504
rect 464 502 466 504
rect 513 502 515 504
rect 557 502 559 504
rect 565 502 567 504
rect 636 502 638 504
rect 35 370 37 372
rect 43 370 45 372
rect 70 370 72 372
rect 119 370 121 372
rect 200 370 202 372
rect 218 370 220 372
rect 230 370 232 372
rect 246 370 248 372
rect 334 370 336 372
rect 448 370 450 372
rect 465 370 467 372
rect 477 370 479 372
rect 521 370 523 372
rect 541 370 543 372
rect 581 370 583 372
rect 122 358 124 360
rect 162 358 164 360
rect 182 358 184 360
rect 226 358 228 360
rect 238 358 240 360
rect 255 358 257 360
rect 369 358 371 360
rect 457 358 459 360
rect 473 358 475 360
rect 485 358 487 360
rect 503 358 505 360
rect 584 358 586 360
rect 633 358 635 360
rect 660 358 662 360
rect 668 358 670 360
rect 67 226 69 228
rect 138 226 140 228
rect 146 226 148 228
rect 190 226 192 228
rect 239 226 241 228
rect 274 226 276 228
rect 286 226 288 228
rect 453 226 455 228
rect 530 226 532 228
rect 605 226 607 228
rect 621 226 623 228
rect 633 226 635 228
rect 84 214 86 216
rect 96 214 98 216
rect 114 214 116 216
rect 493 214 495 216
rect 636 214 638 216
rect 67 82 69 84
rect 168 82 170 84
rect 188 82 190 84
rect 200 82 202 84
rect 429 82 431 84
rect 451 82 453 84
rect 517 82 519 84
rect 605 82 607 84
rect 621 82 623 84
rect 633 82 635 84
rect 82 70 84 72
rect 94 70 96 72
rect 132 70 134 72
rect 184 70 186 72
rect 379 70 381 72
rect 391 70 393 72
rect 488 70 490 72
rect 565 70 567 72
rect 636 70 638 72
<< ptiect1 >>
rect 34 718 36 720
rect 122 718 124 720
rect 138 718 140 720
rect 182 718 184 720
rect 312 718 314 720
rect 324 718 326 720
rect 500 718 502 720
rect 520 718 522 720
rect 538 718 540 720
rect 609 718 611 720
rect 621 718 623 720
rect 633 718 635 720
rect 70 586 72 588
rect 82 586 84 588
rect 98 586 100 588
rect 142 586 144 588
rect 274 586 276 588
rect 503 586 505 588
rect 515 586 517 588
rect 535 586 537 588
rect 669 586 671 588
rect 34 574 36 576
rect 146 574 148 576
rect 254 574 256 576
rect 445 574 447 576
rect 457 574 459 576
rect 509 574 511 576
rect 589 574 591 576
rect 607 574 609 576
rect 619 574 621 576
rect 633 574 635 576
rect 54 442 56 444
rect 70 442 72 444
rect 82 442 84 444
rect 98 442 100 444
rect 206 442 208 444
rect 250 442 252 444
rect 497 442 499 444
rect 513 442 515 444
rect 557 442 559 444
rect 669 442 671 444
rect 70 430 72 432
rect 119 430 121 432
rect 200 430 202 432
rect 218 430 220 432
rect 230 430 232 432
rect 246 430 248 432
rect 290 430 292 432
rect 448 430 450 432
rect 465 430 467 432
rect 477 430 479 432
rect 521 430 523 432
rect 541 430 543 432
rect 625 430 627 432
rect 78 298 80 300
rect 162 298 164 300
rect 182 298 184 300
rect 226 298 228 300
rect 238 298 240 300
rect 255 298 257 300
rect 413 298 415 300
rect 457 298 459 300
rect 473 298 475 300
rect 485 298 487 300
rect 503 298 505 300
rect 584 298 586 300
rect 633 298 635 300
rect 34 286 36 288
rect 146 286 148 288
rect 190 286 192 288
rect 206 286 208 288
rect 274 286 276 288
rect 286 286 288 288
rect 453 286 455 288
rect 497 286 499 288
rect 605 286 607 288
rect 621 286 623 288
rect 633 286 635 288
rect 649 286 651 288
rect 70 154 72 156
rect 84 154 86 156
rect 96 154 98 156
rect 114 154 116 156
rect 194 154 196 156
rect 449 154 451 156
rect 557 154 559 156
rect 669 154 671 156
rect 34 142 36 144
rect 168 142 170 144
rect 188 142 190 144
rect 200 142 202 144
rect 429 142 431 144
rect 561 142 563 144
rect 605 142 607 144
rect 621 142 623 144
rect 633 142 635 144
rect 70 10 72 12
rect 82 10 84 12
rect 94 10 96 12
rect 165 10 167 12
rect 183 10 185 12
rect 203 10 205 12
rect 379 10 381 12
rect 391 10 393 12
rect 521 10 523 12
rect 565 10 567 12
rect 581 10 583 12
rect 669 10 671 12
<< pdifct0 >>
rect 41 682 43 684
rect 51 668 53 670
rect 67 682 69 684
rect 67 675 69 677
rect 51 661 53 663
rect 87 667 89 669
rect 123 668 125 670
rect 189 682 191 684
rect 147 670 149 672
rect 157 675 159 677
rect 157 668 159 670
rect 167 668 169 670
rect 123 661 125 663
rect 199 668 201 670
rect 215 682 217 684
rect 215 675 217 677
rect 199 661 201 663
rect 235 667 237 669
rect 251 665 253 667
rect 261 668 263 670
rect 271 665 273 667
rect 322 668 324 670
rect 500 669 502 671
rect 500 662 502 664
rect 545 682 547 684
rect 520 677 522 679
rect 520 670 522 672
rect 555 668 557 670
rect 571 682 573 684
rect 571 675 573 677
rect 555 661 557 663
rect 591 667 593 669
rect 619 668 621 670
rect 636 668 638 670
rect 636 661 638 663
rect 670 668 672 670
rect 670 661 672 663
rect 33 643 35 645
rect 33 636 35 638
rect 43 636 45 638
rect 43 629 45 631
rect 53 643 55 645
rect 53 636 55 638
rect 80 636 82 638
rect 107 634 109 636
rect 117 636 119 638
rect 117 629 119 631
rect 127 636 129 638
rect 151 635 153 637
rect 161 635 163 637
rect 161 628 163 630
rect 183 634 185 636
rect 183 627 185 629
rect 275 634 277 636
rect 275 627 277 629
rect 505 636 507 638
rect 582 643 584 645
rect 544 634 546 636
rect 554 636 556 638
rect 554 629 556 631
rect 564 636 566 638
rect 582 636 584 638
rect 592 636 594 638
rect 592 629 594 631
rect 602 643 604 645
rect 602 636 604 638
rect 616 637 618 639
rect 652 643 654 645
rect 636 629 638 631
rect 636 622 638 624
rect 652 636 654 638
rect 662 622 664 624
rect 41 538 43 540
rect 51 524 53 526
rect 67 538 69 540
rect 67 531 69 533
rect 51 517 53 519
rect 87 523 89 525
rect 101 524 103 526
rect 101 517 103 519
rect 111 531 113 533
rect 111 524 113 526
rect 121 524 123 526
rect 121 517 123 519
rect 145 524 147 526
rect 145 517 147 519
rect 169 524 171 526
rect 193 524 195 526
rect 213 533 215 535
rect 213 526 215 528
rect 235 532 237 534
rect 235 525 237 527
rect 245 525 247 527
rect 193 517 195 519
rect 455 524 457 526
rect 512 524 514 526
rect 512 517 514 519
rect 546 524 548 526
rect 560 524 562 526
rect 570 531 572 533
rect 570 524 572 526
rect 580 526 582 528
rect 546 517 548 519
rect 617 524 619 526
rect 636 524 638 526
rect 636 517 638 519
rect 670 524 672 526
rect 670 517 672 519
rect 55 499 57 501
rect 55 492 57 494
rect 80 492 82 494
rect 107 490 109 492
rect 117 492 119 494
rect 117 485 119 487
rect 127 492 129 494
rect 153 493 155 495
rect 189 499 191 501
rect 173 485 175 487
rect 173 478 175 480
rect 189 492 191 494
rect 221 492 223 494
rect 231 492 233 494
rect 231 485 233 487
rect 241 490 243 492
rect 199 478 201 480
rect 444 493 446 495
rect 480 499 482 501
rect 464 485 466 487
rect 464 478 466 480
rect 480 492 482 494
rect 490 478 492 480
rect 522 490 524 492
rect 532 492 534 494
rect 532 485 534 487
rect 542 492 544 494
rect 557 490 559 492
rect 577 490 579 492
rect 577 483 579 485
rect 597 490 599 492
rect 616 493 618 495
rect 597 483 599 485
rect 652 499 654 501
rect 636 485 638 487
rect 636 478 638 480
rect 652 492 654 494
rect 662 478 664 480
rect 34 389 36 391
rect 34 382 36 384
rect 45 389 47 391
rect 45 382 47 384
rect 56 380 58 382
rect 79 382 81 384
rect 89 387 91 389
rect 89 380 91 382
rect 99 380 101 382
rect 128 382 130 384
rect 138 387 140 389
rect 138 380 140 382
rect 148 380 150 382
rect 171 380 173 382
rect 181 387 183 389
rect 181 380 183 382
rect 191 382 193 384
rect 228 380 230 382
rect 255 382 257 384
rect 265 387 267 389
rect 265 380 267 382
rect 275 380 277 382
rect 299 381 301 383
rect 309 388 311 390
rect 309 381 311 383
rect 331 389 333 391
rect 331 382 333 384
rect 419 380 421 382
rect 429 387 431 389
rect 429 380 431 382
rect 439 382 441 384
rect 475 380 477 382
rect 492 380 494 382
rect 502 387 504 389
rect 502 380 504 382
rect 512 382 514 384
rect 550 382 552 384
rect 560 387 562 389
rect 560 380 562 382
rect 570 380 572 382
rect 584 389 586 391
rect 584 382 586 384
rect 606 388 608 390
rect 606 381 608 383
rect 616 381 618 383
rect 640 380 642 382
rect 640 373 642 375
rect 660 380 662 382
rect 660 373 662 375
rect 43 355 45 357
rect 43 348 45 350
rect 63 355 65 357
rect 63 348 65 350
rect 87 347 89 349
rect 97 347 99 349
rect 97 340 99 342
rect 119 346 121 348
rect 119 339 121 341
rect 133 348 135 350
rect 143 348 145 350
rect 143 341 145 343
rect 153 346 155 348
rect 191 346 193 348
rect 201 348 203 350
rect 201 341 203 343
rect 211 348 213 350
rect 228 348 230 350
rect 264 346 266 348
rect 274 348 276 350
rect 274 341 276 343
rect 284 348 286 350
rect 372 346 374 348
rect 372 339 374 341
rect 394 347 396 349
rect 394 340 396 342
rect 404 347 406 349
rect 428 348 430 350
rect 438 348 440 350
rect 438 341 440 343
rect 448 346 450 348
rect 475 348 477 350
rect 512 346 514 348
rect 522 348 524 350
rect 522 341 524 343
rect 532 348 534 350
rect 555 348 557 350
rect 565 348 567 350
rect 565 341 567 343
rect 575 346 577 348
rect 604 348 606 350
rect 614 348 616 350
rect 614 341 616 343
rect 624 346 626 348
rect 647 348 649 350
rect 658 346 660 348
rect 658 339 660 341
rect 669 346 671 348
rect 669 339 671 341
rect 41 250 43 252
rect 51 236 53 238
rect 67 250 69 252
rect 67 243 69 245
rect 51 229 53 231
rect 106 245 108 247
rect 87 235 89 237
rect 106 238 108 240
rect 126 245 128 247
rect 126 238 128 240
rect 146 238 148 240
rect 161 236 163 238
rect 171 243 173 245
rect 171 236 173 238
rect 181 238 183 240
rect 213 250 215 252
rect 223 236 225 238
rect 239 250 241 252
rect 239 243 241 245
rect 223 229 225 231
rect 259 235 261 237
rect 284 236 286 238
rect 504 250 506 252
rect 462 238 464 240
rect 472 243 474 245
rect 472 236 474 238
rect 482 236 484 238
rect 514 236 516 238
rect 530 250 532 252
rect 530 243 532 245
rect 514 229 516 231
rect 550 235 552 237
rect 576 236 578 238
rect 586 243 588 245
rect 586 236 588 238
rect 596 238 598 240
rect 623 236 625 238
rect 648 236 650 238
rect 648 229 650 231
rect 33 211 35 213
rect 33 204 35 206
rect 67 211 69 213
rect 67 204 69 206
rect 86 204 88 206
rect 157 211 159 213
rect 123 202 125 204
rect 133 204 135 206
rect 133 197 135 199
rect 143 204 145 206
rect 157 204 159 206
rect 191 211 193 213
rect 510 211 512 213
rect 191 204 193 206
rect 458 203 460 205
rect 468 203 470 205
rect 468 196 470 198
rect 490 202 492 204
rect 490 195 492 197
rect 510 204 512 206
rect 534 204 536 206
rect 558 211 560 213
rect 558 204 560 206
rect 582 211 584 213
rect 582 204 584 206
rect 592 204 594 206
rect 592 197 594 199
rect 602 211 604 213
rect 602 204 604 206
rect 616 205 618 207
rect 652 211 654 213
rect 636 197 638 199
rect 636 190 638 192
rect 652 204 654 206
rect 662 190 664 192
rect 41 106 43 108
rect 51 92 53 94
rect 67 106 69 108
rect 67 99 69 101
rect 51 85 53 87
rect 87 91 89 93
rect 101 92 103 94
rect 101 85 103 87
rect 111 99 113 101
rect 111 92 113 94
rect 121 92 123 94
rect 139 92 141 94
rect 149 99 151 101
rect 149 92 151 94
rect 159 94 161 96
rect 121 85 123 87
rect 198 92 200 94
rect 428 101 430 103
rect 428 94 430 96
rect 520 101 522 103
rect 520 94 522 96
rect 542 100 544 102
rect 542 93 544 95
rect 552 93 554 95
rect 576 92 578 94
rect 586 99 588 101
rect 586 92 588 94
rect 596 94 598 96
rect 623 92 625 94
rect 650 92 652 94
rect 650 85 652 87
rect 660 99 662 101
rect 660 92 662 94
rect 670 92 672 94
rect 670 85 672 87
rect 33 67 35 69
rect 33 60 35 62
rect 67 67 69 69
rect 67 60 69 62
rect 84 60 86 62
rect 112 61 114 63
rect 148 67 150 69
rect 132 53 134 55
rect 132 46 134 48
rect 148 60 150 62
rect 183 58 185 60
rect 183 51 185 53
rect 158 46 160 48
rect 203 66 205 68
rect 203 59 205 61
rect 381 60 383 62
rect 432 63 434 65
rect 442 60 444 62
rect 452 63 454 65
rect 468 61 470 63
rect 504 67 506 69
rect 488 53 490 55
rect 488 46 490 48
rect 504 60 506 62
rect 580 67 582 69
rect 536 60 538 62
rect 546 60 548 62
rect 546 53 548 55
rect 556 58 558 60
rect 514 46 516 48
rect 580 60 582 62
rect 616 61 618 63
rect 652 67 654 69
rect 636 53 638 55
rect 636 46 638 48
rect 652 60 654 62
rect 662 46 664 48
<< pdifct1 >>
rect 77 675 79 677
rect 104 675 106 677
rect 104 668 106 670
rect 137 682 139 684
rect 137 675 139 677
rect 225 675 227 677
rect 311 683 313 685
rect 261 675 263 677
rect 281 675 283 677
rect 281 668 283 670
rect 311 676 313 678
rect 292 658 294 660
rect 510 676 512 678
rect 581 675 583 677
rect 608 683 610 685
rect 608 676 610 678
rect 653 682 655 684
rect 653 675 655 677
rect 172 646 174 648
rect 69 628 71 630
rect 69 621 71 623
rect 97 629 99 631
rect 97 622 99 624
rect 212 646 214 648
rect 141 630 143 632
rect 141 623 143 625
rect 244 628 246 630
rect 516 628 518 630
rect 516 621 518 623
rect 534 629 536 631
rect 534 622 536 624
rect 626 629 628 631
rect 77 531 79 533
rect 169 531 171 533
rect 255 537 257 539
rect 255 530 257 532
rect 444 539 446 541
rect 444 532 446 534
rect 224 514 226 516
rect 529 538 531 540
rect 529 531 531 533
rect 590 538 592 540
rect 590 531 592 533
rect 606 539 608 541
rect 606 532 608 534
rect 653 538 655 540
rect 653 531 655 533
rect 36 492 38 494
rect 36 485 38 487
rect 69 484 71 486
rect 69 477 71 479
rect 97 485 99 487
rect 97 478 99 480
rect 163 485 165 487
rect 251 485 253 487
rect 251 478 253 480
rect 454 485 456 487
rect 512 485 514 487
rect 512 478 514 480
rect 567 485 569 487
rect 567 478 569 480
rect 587 485 589 487
rect 587 478 589 480
rect 626 485 628 487
rect 69 394 71 396
rect 69 387 71 389
rect 118 394 120 396
rect 118 387 120 389
rect 201 394 203 396
rect 201 387 203 389
rect 217 395 219 397
rect 217 388 219 390
rect 245 394 247 396
rect 245 387 247 389
rect 289 393 291 395
rect 289 386 291 388
rect 449 394 451 396
rect 449 387 451 389
rect 464 395 466 397
rect 464 388 466 390
rect 320 370 322 372
rect 522 394 524 396
rect 522 387 524 389
rect 540 394 542 396
rect 540 387 542 389
rect 626 393 628 395
rect 626 386 628 388
rect 595 370 597 372
rect 650 387 652 389
rect 650 380 652 382
rect 670 387 672 389
rect 670 380 672 382
rect 33 348 35 350
rect 33 341 35 343
rect 53 348 55 350
rect 53 341 55 343
rect 108 358 110 360
rect 77 342 79 344
rect 77 335 79 337
rect 163 341 165 343
rect 163 334 165 336
rect 181 341 183 343
rect 181 334 183 336
rect 383 358 385 360
rect 239 340 241 342
rect 239 333 241 335
rect 254 341 256 343
rect 254 334 256 336
rect 414 342 416 344
rect 414 335 416 337
rect 458 341 460 343
rect 458 334 460 336
rect 486 340 488 342
rect 486 333 488 335
rect 502 341 504 343
rect 502 334 504 336
rect 585 341 587 343
rect 585 334 587 336
rect 634 341 636 343
rect 634 334 636 336
rect 77 243 79 245
rect 116 250 118 252
rect 116 243 118 245
rect 136 250 138 252
rect 136 243 138 245
rect 191 250 193 252
rect 191 243 193 245
rect 249 243 251 245
rect 273 251 275 253
rect 273 244 275 246
rect 452 250 454 252
rect 452 243 454 245
rect 540 243 542 245
rect 606 250 608 252
rect 606 243 608 245
rect 634 251 636 253
rect 634 244 636 246
rect 667 243 669 245
rect 667 236 669 238
rect 50 197 52 199
rect 50 190 52 192
rect 97 196 99 198
rect 97 189 99 191
rect 113 197 115 199
rect 113 190 115 192
rect 174 197 176 199
rect 174 190 176 192
rect 479 214 481 216
rect 448 198 450 200
rect 448 191 450 193
rect 534 197 536 199
rect 626 197 628 199
rect 77 99 79 101
rect 169 106 171 108
rect 169 99 171 101
rect 187 107 189 109
rect 187 100 189 102
rect 459 100 461 102
rect 562 105 564 107
rect 562 98 564 100
rect 491 82 493 84
rect 606 106 608 108
rect 606 99 608 101
rect 634 107 636 109
rect 634 100 636 102
rect 531 82 533 84
rect 50 53 52 55
rect 50 46 52 48
rect 95 52 97 54
rect 95 45 97 47
rect 122 53 124 55
rect 193 52 195 54
rect 411 70 413 72
rect 392 52 394 54
rect 422 60 424 62
rect 422 53 424 55
rect 442 53 444 55
rect 392 45 394 47
rect 478 53 480 55
rect 566 53 568 55
rect 566 46 568 48
rect 599 60 601 62
rect 599 53 601 55
rect 626 53 628 55
<< alu0 >>
rect 45 711 51 717
rect 45 709 47 711
rect 49 709 51 711
rect 45 708 51 709
rect 58 708 62 710
rect 58 706 59 708
rect 61 706 62 708
rect 32 703 36 705
rect 32 701 33 703
rect 35 701 36 703
rect 32 695 36 701
rect 58 703 62 706
rect 58 699 82 703
rect 32 691 43 695
rect 39 685 43 691
rect 78 695 82 699
rect 58 694 74 695
rect 58 692 70 694
rect 72 692 74 694
rect 58 691 74 692
rect 78 693 83 695
rect 78 691 80 693
rect 82 691 83 693
rect 58 685 62 691
rect 78 689 83 691
rect 78 687 82 689
rect 39 684 62 685
rect 39 682 41 684
rect 43 682 62 684
rect 39 681 62 682
rect 50 670 54 672
rect 50 668 51 670
rect 53 668 54 670
rect 50 663 54 668
rect 58 670 62 681
rect 66 684 82 687
rect 66 682 67 684
rect 69 683 82 684
rect 69 682 70 683
rect 66 677 70 682
rect 66 675 67 677
rect 69 675 70 677
rect 66 673 70 675
rect 122 708 126 717
rect 122 706 123 708
rect 125 706 126 708
rect 122 704 126 706
rect 193 711 199 717
rect 151 710 171 711
rect 151 708 167 710
rect 169 708 171 710
rect 193 709 195 711
rect 197 709 199 711
rect 193 708 199 709
rect 206 708 210 710
rect 151 707 171 708
rect 139 704 140 706
rect 151 703 155 707
rect 206 706 207 708
rect 209 706 210 708
rect 143 699 155 703
rect 143 694 147 699
rect 143 692 144 694
rect 146 692 147 694
rect 143 680 147 692
rect 180 703 184 705
rect 180 701 181 703
rect 183 701 184 703
rect 180 695 184 701
rect 206 703 210 706
rect 206 699 230 703
rect 180 691 191 695
rect 143 677 160 680
rect 143 676 157 677
rect 156 675 157 676
rect 159 675 160 677
rect 145 672 151 673
rect 58 669 91 670
rect 58 667 87 669
rect 89 667 91 669
rect 122 670 126 672
rect 122 668 123 670
rect 125 668 126 670
rect 58 666 91 667
rect 50 661 51 663
rect 53 661 54 663
rect 122 663 126 668
rect 122 661 123 663
rect 125 661 126 663
rect 145 670 147 672
rect 149 670 151 672
rect 145 661 151 670
rect 156 670 160 675
rect 187 685 191 691
rect 226 695 230 699
rect 206 694 222 695
rect 206 692 218 694
rect 220 692 222 694
rect 206 691 222 692
rect 226 693 231 695
rect 226 691 228 693
rect 230 691 231 693
rect 206 685 210 691
rect 226 689 231 691
rect 226 687 230 689
rect 187 684 210 685
rect 187 682 189 684
rect 191 682 210 684
rect 187 681 210 682
rect 156 668 157 670
rect 159 668 160 670
rect 156 666 160 668
rect 165 670 171 671
rect 165 668 167 670
rect 169 668 171 670
rect 165 661 171 668
rect 198 670 202 672
rect 198 668 199 670
rect 201 668 202 670
rect 198 663 202 668
rect 206 670 210 681
rect 214 684 230 687
rect 214 682 215 684
rect 217 683 230 684
rect 217 682 218 683
rect 214 677 218 682
rect 214 675 215 677
rect 217 675 218 677
rect 214 673 218 675
rect 276 687 281 688
rect 276 685 278 687
rect 280 685 281 687
rect 324 706 328 717
rect 497 710 503 717
rect 497 708 499 710
rect 501 708 503 710
rect 497 707 503 708
rect 520 707 524 717
rect 549 711 555 717
rect 549 709 551 711
rect 553 709 555 711
rect 549 708 555 709
rect 562 708 566 710
rect 276 684 281 685
rect 260 670 264 674
rect 206 669 239 670
rect 206 667 235 669
rect 237 667 239 669
rect 206 666 239 667
rect 250 667 254 669
rect 198 661 199 663
rect 201 661 202 663
rect 250 665 251 667
rect 253 665 254 667
rect 260 668 261 670
rect 263 668 264 670
rect 260 666 264 668
rect 270 667 274 669
rect 250 661 254 665
rect 270 665 271 667
rect 273 665 274 667
rect 313 699 314 705
rect 324 704 325 706
rect 327 704 328 706
rect 520 705 521 707
rect 523 705 524 707
rect 562 706 563 708
rect 565 706 566 708
rect 324 702 328 704
rect 520 703 524 705
rect 536 703 540 705
rect 536 701 537 703
rect 539 701 540 703
rect 313 680 314 687
rect 519 687 521 694
rect 536 695 540 701
rect 562 703 566 706
rect 562 699 586 703
rect 536 691 547 695
rect 518 679 524 680
rect 518 677 520 679
rect 522 677 524 679
rect 518 672 524 677
rect 498 671 504 672
rect 320 670 326 671
rect 320 668 322 670
rect 324 668 326 670
rect 270 661 274 665
rect 320 661 326 668
rect 498 669 500 671
rect 502 669 504 671
rect 498 664 504 669
rect 498 662 500 664
rect 502 662 504 664
rect 498 661 504 662
rect 518 670 520 672
rect 522 670 524 672
rect 518 661 524 670
rect 543 685 547 691
rect 582 695 586 699
rect 562 694 578 695
rect 562 692 574 694
rect 576 692 578 694
rect 562 691 578 692
rect 582 693 587 695
rect 582 691 584 693
rect 586 691 587 693
rect 562 685 566 691
rect 582 689 587 691
rect 582 687 586 689
rect 543 684 566 685
rect 543 682 545 684
rect 547 682 566 684
rect 543 681 566 682
rect 554 670 558 672
rect 554 668 555 670
rect 557 668 558 670
rect 554 663 558 668
rect 562 670 566 681
rect 570 684 586 687
rect 570 682 571 684
rect 573 683 586 684
rect 573 682 574 683
rect 570 677 574 682
rect 570 675 571 677
rect 573 675 574 677
rect 570 673 574 675
rect 621 706 625 717
rect 646 715 648 717
rect 650 715 652 717
rect 610 699 611 705
rect 621 704 622 706
rect 624 704 625 706
rect 621 702 625 704
rect 646 710 652 715
rect 666 715 668 717
rect 670 715 672 717
rect 666 714 672 715
rect 646 708 648 710
rect 650 708 652 710
rect 646 707 652 708
rect 610 680 611 687
rect 617 670 623 671
rect 562 669 595 670
rect 562 667 591 669
rect 593 667 595 669
rect 562 666 595 667
rect 617 668 619 670
rect 621 668 623 670
rect 554 661 555 663
rect 557 661 558 663
rect 617 661 623 668
rect 634 670 640 671
rect 634 668 636 670
rect 638 668 640 670
rect 634 663 640 668
rect 634 661 636 663
rect 638 661 640 663
rect 668 670 674 671
rect 668 668 670 670
rect 672 668 674 670
rect 668 663 674 668
rect 668 661 670 663
rect 672 661 674 663
rect 31 643 33 645
rect 35 643 37 645
rect 31 638 37 643
rect 51 643 53 645
rect 55 643 57 645
rect 31 636 33 638
rect 35 636 37 638
rect 31 635 37 636
rect 42 638 46 640
rect 42 636 43 638
rect 45 636 46 638
rect 42 632 46 636
rect 51 638 57 643
rect 51 636 53 638
rect 55 636 57 638
rect 51 635 57 636
rect 78 638 84 645
rect 78 636 80 638
rect 82 636 84 638
rect 78 635 84 636
rect 105 636 111 645
rect 105 634 107 636
rect 109 634 111 636
rect 105 633 111 634
rect 116 638 120 640
rect 116 636 117 638
rect 119 636 120 638
rect 43 631 46 632
rect 45 629 46 631
rect 43 627 46 629
rect 116 631 120 636
rect 125 638 131 645
rect 125 636 127 638
rect 129 636 131 638
rect 125 635 131 636
rect 149 637 155 645
rect 149 635 151 637
rect 153 635 155 637
rect 149 634 155 635
rect 160 637 187 639
rect 160 635 161 637
rect 163 636 187 637
rect 163 635 183 636
rect 116 630 117 631
rect 54 614 55 618
rect 71 619 72 626
rect 103 629 117 630
rect 119 629 120 631
rect 103 626 120 629
rect 54 598 58 600
rect 54 596 55 598
rect 57 596 58 598
rect 54 591 58 596
rect 71 601 72 607
rect 82 602 86 604
rect 82 600 83 602
rect 85 600 86 602
rect 54 589 55 591
rect 57 589 58 591
rect 82 589 86 600
rect 103 614 107 626
rect 160 630 164 635
rect 181 634 183 635
rect 185 634 187 636
rect 155 628 161 630
rect 163 628 164 630
rect 103 612 104 614
rect 106 612 107 614
rect 103 607 107 612
rect 103 603 115 607
rect 99 600 100 602
rect 111 599 115 603
rect 143 621 144 627
rect 155 626 164 628
rect 155 623 159 626
rect 181 629 187 634
rect 181 627 183 629
rect 185 627 187 629
rect 181 626 187 627
rect 147 619 159 623
rect 147 614 151 619
rect 166 618 172 619
rect 147 612 148 614
rect 150 612 151 614
rect 147 606 151 612
rect 111 598 131 599
rect 111 596 127 598
rect 129 596 131 598
rect 111 595 131 596
rect 143 600 144 606
rect 147 602 156 606
rect 211 611 212 617
rect 152 598 156 602
rect 273 636 279 645
rect 273 634 275 636
rect 277 634 279 636
rect 503 638 509 645
rect 503 636 505 638
rect 507 636 509 638
rect 503 635 509 636
rect 542 636 548 645
rect 273 629 279 634
rect 542 634 544 636
rect 546 634 548 636
rect 542 633 548 634
rect 553 638 557 640
rect 553 636 554 638
rect 556 636 557 638
rect 273 627 275 629
rect 277 627 279 629
rect 273 626 279 627
rect 515 619 516 626
rect 152 597 182 598
rect 152 595 178 597
rect 180 595 182 597
rect 152 594 182 595
rect 208 597 212 599
rect 208 595 209 597
rect 211 595 212 597
rect 208 589 212 595
rect 250 597 254 599
rect 250 595 251 597
rect 253 595 254 597
rect 250 589 254 595
rect 501 602 505 604
rect 501 600 502 602
rect 504 600 505 602
rect 515 601 516 607
rect 501 589 505 600
rect 553 631 557 636
rect 562 638 568 645
rect 562 636 564 638
rect 566 636 568 638
rect 562 635 568 636
rect 580 643 582 645
rect 584 643 586 645
rect 580 638 586 643
rect 600 643 602 645
rect 604 643 606 645
rect 580 636 582 638
rect 584 636 586 638
rect 580 635 586 636
rect 591 638 595 640
rect 591 636 592 638
rect 594 636 595 638
rect 591 632 595 636
rect 600 638 606 643
rect 651 643 652 645
rect 654 643 655 645
rect 600 636 602 638
rect 604 636 606 638
rect 614 639 647 640
rect 614 637 616 639
rect 618 637 647 639
rect 614 636 647 637
rect 600 635 606 636
rect 553 630 554 631
rect 540 629 554 630
rect 556 629 557 631
rect 540 626 557 629
rect 540 614 544 626
rect 591 631 594 632
rect 591 629 592 631
rect 591 627 594 629
rect 540 612 541 614
rect 543 612 544 614
rect 540 607 544 612
rect 540 603 552 607
rect 536 600 537 602
rect 548 599 552 603
rect 582 614 583 618
rect 548 598 568 599
rect 548 596 564 598
rect 566 596 568 598
rect 548 595 568 596
rect 579 598 583 600
rect 579 596 580 598
rect 582 596 583 598
rect 579 591 583 596
rect 635 631 639 633
rect 635 629 636 631
rect 638 629 639 631
rect 635 624 639 629
rect 635 623 636 624
rect 623 622 636 623
rect 638 622 639 624
rect 623 619 639 622
rect 643 625 647 636
rect 651 638 655 643
rect 651 636 652 638
rect 654 636 655 638
rect 651 634 655 636
rect 643 624 666 625
rect 643 622 662 624
rect 664 622 666 624
rect 643 621 666 622
rect 623 617 627 619
rect 622 615 627 617
rect 643 615 647 621
rect 622 613 623 615
rect 625 613 627 615
rect 622 611 627 613
rect 631 614 647 615
rect 631 612 633 614
rect 635 612 647 614
rect 631 611 647 612
rect 623 607 627 611
rect 662 615 666 621
rect 662 611 673 615
rect 623 603 647 607
rect 643 600 647 603
rect 669 605 673 611
rect 669 603 670 605
rect 672 603 673 605
rect 669 601 673 603
rect 643 598 644 600
rect 646 598 647 600
rect 643 596 647 598
rect 654 597 660 598
rect 654 595 656 597
rect 658 595 660 597
rect 579 589 580 591
rect 582 589 583 591
rect 654 589 660 595
rect 45 567 51 573
rect 122 571 123 573
rect 125 571 126 573
rect 45 565 47 567
rect 49 565 51 567
rect 45 564 51 565
rect 58 564 62 566
rect 58 562 59 564
rect 61 562 62 564
rect 32 559 36 561
rect 32 557 33 559
rect 35 557 36 559
rect 32 551 36 557
rect 58 559 62 562
rect 58 555 82 559
rect 32 547 43 551
rect 39 541 43 547
rect 78 551 82 555
rect 58 550 74 551
rect 58 548 70 550
rect 72 548 74 550
rect 58 547 74 548
rect 78 549 83 551
rect 78 547 80 549
rect 82 547 83 549
rect 58 541 62 547
rect 78 545 83 547
rect 78 543 82 545
rect 39 540 62 541
rect 39 538 41 540
rect 43 538 62 540
rect 39 537 62 538
rect 50 526 54 528
rect 50 524 51 526
rect 53 524 54 526
rect 50 519 54 524
rect 58 526 62 537
rect 66 540 82 543
rect 66 538 67 540
rect 69 539 82 540
rect 69 538 70 539
rect 66 533 70 538
rect 66 531 67 533
rect 69 531 70 533
rect 66 529 70 531
rect 122 566 126 571
rect 122 564 123 566
rect 125 564 126 566
rect 122 562 126 564
rect 216 567 246 568
rect 216 565 218 567
rect 220 565 246 567
rect 216 564 246 565
rect 122 544 123 548
rect 242 560 246 564
rect 242 556 251 560
rect 254 556 255 562
rect 247 550 251 556
rect 247 548 248 550
rect 250 548 251 550
rect 226 543 232 544
rect 247 543 251 548
rect 239 539 251 543
rect 111 533 114 535
rect 113 531 114 533
rect 211 535 217 536
rect 211 533 213 535
rect 215 533 217 535
rect 111 530 114 531
rect 99 526 105 527
rect 58 525 91 526
rect 58 523 87 525
rect 89 523 91 525
rect 58 522 91 523
rect 99 524 101 526
rect 103 524 105 526
rect 50 517 51 519
rect 53 517 54 519
rect 99 519 105 524
rect 110 526 114 530
rect 110 524 111 526
rect 113 524 114 526
rect 110 522 114 524
rect 119 526 125 527
rect 119 524 121 526
rect 123 524 125 526
rect 99 517 101 519
rect 103 517 105 519
rect 119 519 125 524
rect 119 517 121 519
rect 123 517 125 519
rect 143 526 149 527
rect 143 524 145 526
rect 147 524 149 526
rect 143 519 149 524
rect 168 526 172 531
rect 211 528 217 533
rect 239 536 243 539
rect 234 534 243 536
rect 254 535 255 541
rect 234 532 235 534
rect 237 532 243 534
rect 168 524 169 526
rect 171 524 172 526
rect 168 522 172 524
rect 191 526 197 527
rect 191 524 193 526
rect 195 524 197 526
rect 143 517 145 519
rect 147 517 149 519
rect 191 519 197 524
rect 211 526 213 528
rect 215 527 217 528
rect 234 527 238 532
rect 457 562 461 573
rect 522 571 524 573
rect 526 571 528 573
rect 446 555 447 561
rect 457 560 458 562
rect 460 560 461 562
rect 457 558 461 560
rect 522 566 528 571
rect 542 571 544 573
rect 546 571 548 573
rect 542 570 548 571
rect 522 564 524 566
rect 526 564 528 566
rect 522 563 528 564
rect 558 566 578 567
rect 558 564 560 566
rect 562 564 578 566
rect 558 563 578 564
rect 446 536 447 543
rect 574 559 578 563
rect 589 560 590 562
rect 574 555 586 559
rect 582 550 586 555
rect 582 548 583 550
rect 585 548 586 550
rect 215 526 235 527
rect 211 525 235 526
rect 237 525 238 527
rect 211 523 238 525
rect 243 527 249 528
rect 243 525 245 527
rect 247 525 249 527
rect 191 517 193 519
rect 195 517 197 519
rect 243 517 249 525
rect 582 536 586 548
rect 569 533 586 536
rect 569 531 570 533
rect 572 532 586 533
rect 619 562 623 573
rect 646 571 648 573
rect 650 571 652 573
rect 608 555 609 561
rect 619 560 620 562
rect 622 560 623 562
rect 619 558 623 560
rect 646 566 652 571
rect 666 571 668 573
rect 670 571 672 573
rect 666 570 672 571
rect 646 564 648 566
rect 650 564 652 566
rect 646 563 652 564
rect 608 536 609 543
rect 572 531 573 532
rect 453 526 459 527
rect 453 524 455 526
rect 457 524 459 526
rect 453 517 459 524
rect 510 526 516 527
rect 510 524 512 526
rect 514 524 516 526
rect 510 519 516 524
rect 510 517 512 519
rect 514 517 516 519
rect 544 526 550 527
rect 544 524 546 526
rect 548 524 550 526
rect 544 519 550 524
rect 544 517 546 519
rect 548 517 550 519
rect 558 526 564 527
rect 558 524 560 526
rect 562 524 564 526
rect 558 517 564 524
rect 569 526 573 531
rect 569 524 570 526
rect 572 524 573 526
rect 569 522 573 524
rect 578 528 584 529
rect 578 526 580 528
rect 582 526 584 528
rect 578 517 584 526
rect 615 526 621 527
rect 615 524 617 526
rect 619 524 621 526
rect 615 517 621 524
rect 634 526 640 527
rect 634 524 636 526
rect 638 524 640 526
rect 634 519 640 524
rect 634 517 636 519
rect 638 517 640 519
rect 668 526 674 527
rect 668 524 670 526
rect 672 524 674 526
rect 668 519 674 524
rect 668 517 670 519
rect 672 517 674 519
rect 54 499 55 501
rect 57 499 58 501
rect 54 494 58 499
rect 54 492 55 494
rect 57 492 58 494
rect 54 490 58 492
rect 78 494 84 501
rect 78 492 80 494
rect 82 492 84 494
rect 78 491 84 492
rect 105 492 111 501
rect 105 490 107 492
rect 109 490 111 492
rect 105 489 111 490
rect 116 494 120 496
rect 116 492 117 494
rect 119 492 120 494
rect 116 487 120 492
rect 125 494 131 501
rect 188 499 189 501
rect 191 499 192 501
rect 125 492 127 494
rect 129 492 131 494
rect 151 495 184 496
rect 151 493 153 495
rect 155 493 184 495
rect 151 492 184 493
rect 125 491 131 492
rect 116 486 117 487
rect 71 475 72 482
rect 103 485 117 486
rect 119 485 120 487
rect 103 482 120 485
rect 54 456 58 458
rect 54 454 55 456
rect 57 454 58 456
rect 54 445 58 454
rect 71 457 72 463
rect 82 458 86 460
rect 82 456 83 458
rect 85 456 86 458
rect 82 445 86 456
rect 103 470 107 482
rect 172 487 176 489
rect 172 485 173 487
rect 175 485 176 487
rect 103 468 104 470
rect 106 468 107 470
rect 103 463 107 468
rect 103 459 115 463
rect 99 456 100 458
rect 111 455 115 459
rect 111 454 131 455
rect 111 452 127 454
rect 129 452 131 454
rect 111 451 131 452
rect 172 480 176 485
rect 172 479 173 480
rect 160 478 173 479
rect 175 478 176 480
rect 160 475 176 478
rect 180 481 184 492
rect 188 494 192 499
rect 188 492 189 494
rect 191 492 192 494
rect 188 490 192 492
rect 219 494 225 501
rect 219 492 221 494
rect 223 492 225 494
rect 219 491 225 492
rect 230 494 234 496
rect 230 492 231 494
rect 233 492 234 494
rect 180 480 203 481
rect 180 478 199 480
rect 201 478 203 480
rect 180 477 203 478
rect 160 473 164 475
rect 159 471 164 473
rect 180 471 184 477
rect 159 469 160 471
rect 162 469 164 471
rect 159 467 164 469
rect 168 470 184 471
rect 168 468 170 470
rect 172 468 184 470
rect 168 467 184 468
rect 160 463 164 467
rect 199 471 203 477
rect 230 487 234 492
rect 239 492 245 501
rect 479 499 480 501
rect 482 499 483 501
rect 442 495 475 496
rect 442 493 444 495
rect 446 493 475 495
rect 442 492 475 493
rect 239 490 241 492
rect 243 490 245 492
rect 239 489 245 490
rect 230 485 231 487
rect 233 486 234 487
rect 233 485 247 486
rect 230 482 247 485
rect 199 467 210 471
rect 160 459 184 463
rect 180 456 184 459
rect 206 461 210 467
rect 206 459 207 461
rect 209 459 210 461
rect 206 457 210 459
rect 243 470 247 482
rect 243 468 244 470
rect 246 468 247 470
rect 243 463 247 468
rect 235 459 247 463
rect 180 454 181 456
rect 183 454 184 456
rect 235 455 239 459
rect 250 456 251 458
rect 219 454 239 455
rect 180 452 184 454
rect 191 453 197 454
rect 191 451 193 453
rect 195 451 197 453
rect 219 452 221 454
rect 223 452 239 454
rect 219 451 239 452
rect 191 445 197 451
rect 463 487 467 489
rect 463 485 464 487
rect 466 485 467 487
rect 463 480 467 485
rect 463 479 464 480
rect 451 478 464 479
rect 466 478 467 480
rect 451 475 467 478
rect 471 481 475 492
rect 479 494 483 499
rect 479 492 480 494
rect 482 492 483 494
rect 479 490 483 492
rect 471 480 494 481
rect 471 478 490 480
rect 492 478 494 480
rect 471 477 494 478
rect 451 473 455 475
rect 450 471 455 473
rect 471 471 475 477
rect 450 469 451 471
rect 453 469 455 471
rect 450 467 455 469
rect 459 470 475 471
rect 459 468 461 470
rect 463 468 475 470
rect 459 467 475 468
rect 451 463 455 467
rect 490 471 494 477
rect 520 492 526 501
rect 520 490 522 492
rect 524 490 526 492
rect 520 489 526 490
rect 531 494 535 496
rect 531 492 532 494
rect 534 492 535 494
rect 531 487 535 492
rect 540 494 546 501
rect 540 492 542 494
rect 544 492 546 494
rect 540 491 546 492
rect 556 492 560 501
rect 556 490 557 492
rect 559 490 560 492
rect 556 488 560 490
rect 575 492 581 501
rect 575 490 577 492
rect 579 490 581 492
rect 531 486 532 487
rect 518 485 532 486
rect 534 485 535 487
rect 518 482 535 485
rect 490 467 501 471
rect 451 459 475 463
rect 471 456 475 459
rect 497 461 501 467
rect 497 459 498 461
rect 500 459 501 461
rect 497 457 501 459
rect 471 454 472 456
rect 474 454 475 456
rect 518 470 522 482
rect 575 485 581 490
rect 596 492 600 501
rect 651 499 652 501
rect 654 499 655 501
rect 614 495 647 496
rect 614 493 616 495
rect 618 493 647 495
rect 614 492 647 493
rect 596 490 597 492
rect 599 490 600 492
rect 575 483 577 485
rect 579 483 581 485
rect 575 482 581 483
rect 596 485 600 490
rect 596 483 597 485
rect 599 483 600 485
rect 596 481 600 483
rect 635 487 639 489
rect 635 485 636 487
rect 638 485 639 487
rect 518 468 519 470
rect 521 468 522 470
rect 518 463 522 468
rect 518 459 530 463
rect 514 456 515 458
rect 471 452 475 454
rect 482 453 488 454
rect 482 451 484 453
rect 486 451 488 453
rect 482 445 488 451
rect 526 455 530 459
rect 554 461 580 462
rect 554 459 556 461
rect 558 460 580 461
rect 558 459 577 460
rect 554 458 577 459
rect 579 458 580 460
rect 526 454 546 455
rect 575 454 580 458
rect 635 480 639 485
rect 635 479 636 480
rect 623 478 636 479
rect 638 478 639 480
rect 623 475 639 478
rect 643 481 647 492
rect 651 494 655 499
rect 651 492 652 494
rect 654 492 655 494
rect 651 490 655 492
rect 643 480 666 481
rect 643 478 662 480
rect 664 478 666 480
rect 643 477 666 478
rect 623 473 627 475
rect 622 471 627 473
rect 643 471 647 477
rect 622 469 623 471
rect 625 469 627 471
rect 622 467 627 469
rect 631 470 647 471
rect 631 468 633 470
rect 635 468 647 470
rect 631 467 647 468
rect 623 463 627 467
rect 662 471 666 477
rect 662 467 673 471
rect 623 459 647 463
rect 643 456 647 459
rect 669 461 673 467
rect 669 459 670 461
rect 672 459 673 461
rect 669 457 673 459
rect 526 452 542 454
rect 544 452 546 454
rect 526 451 546 452
rect 566 452 570 454
rect 566 450 567 452
rect 569 450 570 452
rect 575 453 601 454
rect 575 451 577 453
rect 579 451 597 453
rect 599 451 601 453
rect 643 454 644 456
rect 646 454 647 456
rect 643 452 647 454
rect 654 453 660 454
rect 654 451 656 453
rect 658 451 660 453
rect 575 450 601 451
rect 566 445 570 450
rect 654 445 660 451
rect 33 428 37 429
rect 33 426 34 428
rect 36 426 37 428
rect 33 424 37 426
rect 32 391 38 392
rect 32 389 34 391
rect 36 389 38 391
rect 32 384 38 389
rect 32 382 34 384
rect 36 382 38 384
rect 32 373 38 382
rect 43 391 56 392
rect 43 389 45 391
rect 43 387 47 389
rect 83 422 103 423
rect 83 420 99 422
rect 101 420 103 422
rect 83 419 103 420
rect 71 416 72 418
rect 83 415 87 419
rect 132 422 152 423
rect 132 420 148 422
rect 150 420 152 422
rect 132 419 152 420
rect 169 422 189 423
rect 169 420 171 422
rect 173 420 189 422
rect 169 419 189 420
rect 75 411 87 415
rect 75 406 79 411
rect 75 404 76 406
rect 78 404 79 406
rect 75 392 79 404
rect 75 389 92 392
rect 75 388 89 389
rect 43 384 49 387
rect 43 382 45 384
rect 47 382 49 384
rect 88 387 89 388
rect 91 387 92 389
rect 43 381 49 382
rect 54 382 60 383
rect 54 380 56 382
rect 58 380 60 382
rect 77 384 83 385
rect 77 382 79 384
rect 81 382 83 384
rect 54 373 60 380
rect 77 373 83 382
rect 88 382 92 387
rect 120 416 121 418
rect 132 415 136 419
rect 124 411 136 415
rect 124 406 128 411
rect 124 404 125 406
rect 127 404 128 406
rect 124 392 128 404
rect 185 415 189 419
rect 200 416 201 418
rect 185 411 197 415
rect 193 406 197 411
rect 193 404 194 406
rect 196 404 197 406
rect 124 389 141 392
rect 124 388 138 389
rect 137 387 138 388
rect 140 387 141 389
rect 126 384 132 385
rect 88 380 89 382
rect 91 380 92 382
rect 88 378 92 380
rect 97 382 103 383
rect 97 380 99 382
rect 101 380 103 382
rect 97 373 103 380
rect 126 382 128 384
rect 130 382 132 384
rect 126 373 132 382
rect 137 382 141 387
rect 193 392 197 404
rect 180 389 197 392
rect 180 387 181 389
rect 183 388 197 389
rect 183 387 184 388
rect 137 380 138 382
rect 140 380 141 382
rect 137 378 141 380
rect 146 382 152 383
rect 146 380 148 382
rect 150 380 152 382
rect 146 373 152 380
rect 169 382 175 383
rect 169 380 171 382
rect 173 380 175 382
rect 169 373 175 380
rect 180 382 184 387
rect 230 418 234 429
rect 219 411 220 417
rect 230 416 231 418
rect 233 416 234 418
rect 230 414 234 416
rect 259 422 279 423
rect 259 420 275 422
rect 277 420 279 422
rect 259 419 279 420
rect 219 392 220 399
rect 247 416 248 418
rect 259 415 263 419
rect 300 423 330 424
rect 300 421 326 423
rect 328 421 330 423
rect 300 420 330 421
rect 417 422 437 423
rect 417 420 419 422
rect 421 420 437 422
rect 251 411 263 415
rect 251 406 255 411
rect 251 404 252 406
rect 254 404 255 406
rect 251 392 255 404
rect 251 389 268 392
rect 251 388 265 389
rect 264 387 265 388
rect 267 387 268 389
rect 180 380 181 382
rect 183 380 184 382
rect 180 378 184 380
rect 189 384 195 385
rect 189 382 191 384
rect 193 382 195 384
rect 253 384 259 385
rect 189 373 195 382
rect 226 382 232 383
rect 226 380 228 382
rect 230 380 232 382
rect 226 373 232 380
rect 253 382 255 384
rect 257 382 259 384
rect 253 373 259 382
rect 264 382 268 387
rect 291 412 292 418
rect 300 416 304 420
rect 417 419 437 420
rect 295 412 304 416
rect 295 406 299 412
rect 295 404 296 406
rect 298 404 299 406
rect 295 399 299 404
rect 433 415 437 419
rect 448 416 449 418
rect 433 411 445 415
rect 441 406 445 411
rect 441 404 442 406
rect 444 404 445 406
rect 314 399 320 400
rect 291 391 292 397
rect 295 395 307 399
rect 303 392 307 395
rect 303 390 312 392
rect 303 388 309 390
rect 311 388 312 390
rect 264 380 265 382
rect 267 380 268 382
rect 264 378 268 380
rect 273 382 279 383
rect 273 380 275 382
rect 277 380 279 382
rect 273 373 279 380
rect 297 383 303 384
rect 297 381 299 383
rect 301 381 303 383
rect 297 373 303 381
rect 308 383 312 388
rect 329 391 335 392
rect 329 389 331 391
rect 333 389 335 391
rect 329 384 335 389
rect 441 392 445 404
rect 428 389 445 392
rect 428 387 429 389
rect 431 388 445 389
rect 431 387 432 388
rect 329 383 331 384
rect 308 381 309 383
rect 311 382 331 383
rect 333 382 335 384
rect 311 381 335 382
rect 308 379 335 381
rect 417 382 423 383
rect 417 380 419 382
rect 421 380 423 382
rect 417 373 423 380
rect 428 382 432 387
rect 477 418 481 429
rect 640 428 642 429
rect 644 428 646 429
rect 640 427 646 428
rect 490 422 510 423
rect 490 420 492 422
rect 494 420 510 422
rect 490 419 510 420
rect 466 411 467 417
rect 477 416 478 418
rect 480 416 481 418
rect 477 414 481 416
rect 506 415 510 419
rect 521 416 522 418
rect 506 411 518 415
rect 514 406 518 411
rect 514 404 515 406
rect 517 404 518 406
rect 466 392 467 399
rect 514 392 518 404
rect 501 389 518 392
rect 501 387 502 389
rect 504 388 518 389
rect 504 387 505 388
rect 428 380 429 382
rect 431 380 432 382
rect 428 378 432 380
rect 437 384 443 385
rect 437 382 439 384
rect 441 382 443 384
rect 437 373 443 382
rect 473 382 479 383
rect 473 380 475 382
rect 477 380 479 382
rect 473 373 479 380
rect 490 382 496 383
rect 490 380 492 382
rect 494 380 496 382
rect 490 373 496 380
rect 501 382 505 387
rect 587 423 617 424
rect 554 422 574 423
rect 554 420 570 422
rect 572 420 574 422
rect 587 421 589 423
rect 591 421 617 423
rect 587 420 617 421
rect 554 419 574 420
rect 542 416 543 418
rect 554 415 558 419
rect 613 416 617 420
rect 546 411 558 415
rect 546 406 550 411
rect 546 404 547 406
rect 549 404 550 406
rect 546 392 550 404
rect 613 412 622 416
rect 625 412 626 418
rect 618 406 622 412
rect 618 404 619 406
rect 621 404 622 406
rect 597 399 603 400
rect 618 399 622 404
rect 610 395 622 399
rect 546 389 563 392
rect 546 388 560 389
rect 559 387 560 388
rect 562 387 563 389
rect 501 380 502 382
rect 504 380 505 382
rect 501 378 505 380
rect 510 384 516 385
rect 510 382 512 384
rect 514 382 516 384
rect 510 373 516 382
rect 548 384 554 385
rect 548 382 550 384
rect 552 382 554 384
rect 548 373 554 382
rect 559 382 563 387
rect 582 391 588 392
rect 582 389 584 391
rect 586 389 588 391
rect 582 384 588 389
rect 610 392 614 395
rect 605 390 614 392
rect 625 391 626 397
rect 605 388 606 390
rect 608 388 614 390
rect 559 380 560 382
rect 562 380 563 382
rect 559 378 563 380
rect 568 382 574 383
rect 568 380 570 382
rect 572 380 574 382
rect 568 373 574 380
rect 582 382 584 384
rect 586 383 588 384
rect 605 383 609 388
rect 586 382 606 383
rect 582 381 606 382
rect 608 381 609 383
rect 582 379 609 381
rect 614 383 620 384
rect 614 381 616 383
rect 618 381 620 383
rect 614 373 620 381
rect 638 382 644 383
rect 638 380 640 382
rect 642 380 644 382
rect 638 375 644 380
rect 658 382 664 383
rect 658 380 660 382
rect 662 380 664 382
rect 638 373 640 375
rect 642 373 644 375
rect 658 375 664 380
rect 658 373 660 375
rect 662 373 664 375
rect 41 355 43 357
rect 45 355 47 357
rect 41 350 47 355
rect 61 355 63 357
rect 65 355 67 357
rect 41 348 43 350
rect 45 348 47 350
rect 41 347 47 348
rect 61 350 67 355
rect 61 348 63 350
rect 65 348 67 350
rect 61 347 67 348
rect 85 349 91 357
rect 85 347 87 349
rect 89 347 91 349
rect 85 346 91 347
rect 96 349 123 351
rect 96 347 97 349
rect 99 348 123 349
rect 99 347 119 348
rect 96 342 100 347
rect 117 346 119 347
rect 121 346 123 348
rect 131 350 137 357
rect 131 348 133 350
rect 135 348 137 350
rect 131 347 137 348
rect 142 350 146 352
rect 142 348 143 350
rect 145 348 146 350
rect 91 340 97 342
rect 99 340 100 342
rect 79 333 80 339
rect 91 338 100 340
rect 91 335 95 338
rect 117 341 123 346
rect 117 339 119 341
rect 121 339 123 341
rect 117 338 123 339
rect 142 343 146 348
rect 151 348 157 357
rect 151 346 153 348
rect 155 346 157 348
rect 151 345 157 346
rect 189 348 195 357
rect 189 346 191 348
rect 193 346 195 348
rect 189 345 195 346
rect 200 350 204 352
rect 200 348 201 350
rect 203 348 204 350
rect 142 341 143 343
rect 145 342 146 343
rect 145 341 159 342
rect 142 338 159 341
rect 83 331 95 335
rect 83 326 87 331
rect 102 330 108 331
rect 83 324 84 326
rect 86 324 87 326
rect 83 318 87 324
rect 79 312 80 318
rect 83 314 92 318
rect 155 326 159 338
rect 155 324 156 326
rect 158 324 159 326
rect 155 319 159 324
rect 147 315 159 319
rect 88 310 92 314
rect 147 311 151 315
rect 162 312 163 314
rect 131 310 151 311
rect 88 309 118 310
rect 88 307 114 309
rect 116 307 118 309
rect 131 308 133 310
rect 135 308 151 310
rect 131 307 151 308
rect 88 306 118 307
rect 200 343 204 348
rect 209 350 215 357
rect 209 348 211 350
rect 213 348 215 350
rect 209 347 215 348
rect 226 350 232 357
rect 226 348 228 350
rect 230 348 232 350
rect 226 347 232 348
rect 262 348 268 357
rect 262 346 264 348
rect 266 346 268 348
rect 262 345 268 346
rect 273 350 277 352
rect 273 348 274 350
rect 276 348 277 350
rect 200 342 201 343
rect 187 341 201 342
rect 203 341 204 343
rect 187 338 204 341
rect 187 326 191 338
rect 238 331 239 338
rect 187 324 188 326
rect 190 324 191 326
rect 187 319 191 324
rect 187 315 199 319
rect 183 312 184 314
rect 195 311 199 315
rect 224 314 228 316
rect 224 312 225 314
rect 227 312 228 314
rect 238 313 239 319
rect 195 310 215 311
rect 195 308 211 310
rect 213 308 215 310
rect 195 307 215 308
rect 59 302 65 303
rect 59 301 61 302
rect 63 301 65 302
rect 224 301 228 312
rect 273 343 277 348
rect 282 350 288 357
rect 282 348 284 350
rect 286 348 288 350
rect 282 347 288 348
rect 370 349 397 351
rect 370 348 394 349
rect 370 346 372 348
rect 374 347 394 348
rect 396 347 397 349
rect 374 346 376 347
rect 273 342 274 343
rect 260 341 274 342
rect 276 341 277 343
rect 260 338 277 341
rect 260 326 264 338
rect 370 341 376 346
rect 370 339 372 341
rect 374 339 376 341
rect 370 338 376 339
rect 393 342 397 347
rect 402 349 408 357
rect 402 347 404 349
rect 406 347 408 349
rect 402 346 408 347
rect 426 350 432 357
rect 426 348 428 350
rect 430 348 432 350
rect 426 347 432 348
rect 437 350 441 352
rect 437 348 438 350
rect 440 348 441 350
rect 393 340 394 342
rect 396 340 402 342
rect 393 338 402 340
rect 398 335 402 338
rect 398 331 410 335
rect 413 333 414 339
rect 385 330 391 331
rect 260 324 261 326
rect 263 324 264 326
rect 260 319 264 324
rect 260 315 272 319
rect 256 312 257 314
rect 268 311 272 315
rect 406 326 410 331
rect 406 324 407 326
rect 409 324 410 326
rect 406 318 410 324
rect 401 314 410 318
rect 268 310 288 311
rect 401 310 405 314
rect 413 312 414 318
rect 437 343 441 348
rect 446 348 452 357
rect 446 346 448 348
rect 450 346 452 348
rect 473 350 479 357
rect 473 348 475 350
rect 477 348 479 350
rect 473 347 479 348
rect 510 348 516 357
rect 446 345 452 346
rect 510 346 512 348
rect 514 346 516 348
rect 510 345 516 346
rect 521 350 525 352
rect 521 348 522 350
rect 524 348 525 350
rect 437 341 438 343
rect 440 342 441 343
rect 440 341 454 342
rect 437 338 454 341
rect 450 326 454 338
rect 450 324 451 326
rect 453 324 454 326
rect 450 319 454 324
rect 442 315 454 319
rect 268 308 284 310
rect 286 308 288 310
rect 268 307 288 308
rect 375 309 405 310
rect 375 307 377 309
rect 379 307 405 309
rect 375 306 405 307
rect 442 311 446 315
rect 457 312 458 314
rect 485 331 486 338
rect 426 310 446 311
rect 426 308 428 310
rect 430 308 446 310
rect 426 307 446 308
rect 471 314 475 316
rect 471 312 472 314
rect 474 312 475 314
rect 485 313 486 319
rect 471 301 475 312
rect 521 343 525 348
rect 530 350 536 357
rect 530 348 532 350
rect 534 348 536 350
rect 530 347 536 348
rect 553 350 559 357
rect 553 348 555 350
rect 557 348 559 350
rect 553 347 559 348
rect 564 350 568 352
rect 564 348 565 350
rect 567 348 568 350
rect 521 342 522 343
rect 508 341 522 342
rect 524 341 525 343
rect 508 338 525 341
rect 508 326 512 338
rect 564 343 568 348
rect 573 348 579 357
rect 573 346 575 348
rect 577 346 579 348
rect 602 350 608 357
rect 602 348 604 350
rect 606 348 608 350
rect 602 347 608 348
rect 613 350 617 352
rect 613 348 614 350
rect 616 348 617 350
rect 573 345 579 346
rect 564 341 565 343
rect 567 342 568 343
rect 567 341 581 342
rect 564 338 581 341
rect 508 324 509 326
rect 511 324 512 326
rect 508 319 512 324
rect 508 315 520 319
rect 504 312 505 314
rect 516 311 520 315
rect 577 326 581 338
rect 577 324 578 326
rect 580 324 581 326
rect 577 319 581 324
rect 569 315 581 319
rect 569 311 573 315
rect 584 312 585 314
rect 613 343 617 348
rect 622 348 628 357
rect 645 350 651 357
rect 622 346 624 348
rect 626 346 628 348
rect 622 345 628 346
rect 645 348 647 350
rect 649 348 651 350
rect 645 347 651 348
rect 656 348 662 349
rect 613 341 614 343
rect 616 342 617 343
rect 656 346 658 348
rect 660 346 662 348
rect 656 343 662 346
rect 616 341 630 342
rect 613 338 630 341
rect 626 326 630 338
rect 626 324 627 326
rect 629 324 630 326
rect 626 319 630 324
rect 618 315 630 319
rect 516 310 536 311
rect 516 308 532 310
rect 534 308 536 310
rect 516 307 536 308
rect 553 310 573 311
rect 553 308 555 310
rect 557 308 573 310
rect 553 307 573 308
rect 618 311 622 315
rect 633 312 634 314
rect 602 310 622 311
rect 602 308 604 310
rect 606 308 622 310
rect 602 307 622 308
rect 658 341 662 343
rect 660 339 662 341
rect 649 338 662 339
rect 667 348 673 357
rect 667 346 669 348
rect 671 346 673 348
rect 667 341 673 346
rect 667 339 669 341
rect 671 339 673 341
rect 667 338 673 339
rect 668 304 672 306
rect 668 302 669 304
rect 671 302 672 304
rect 668 301 672 302
rect 45 279 51 285
rect 135 280 139 285
rect 104 279 130 280
rect 45 277 47 279
rect 49 277 51 279
rect 45 276 51 277
rect 58 276 62 278
rect 58 274 59 276
rect 61 274 62 276
rect 104 277 106 279
rect 108 277 126 279
rect 128 277 130 279
rect 104 276 130 277
rect 135 278 136 280
rect 138 278 139 280
rect 135 276 139 278
rect 159 278 179 279
rect 159 276 161 278
rect 163 276 179 278
rect 32 271 36 273
rect 32 269 33 271
rect 35 269 36 271
rect 32 263 36 269
rect 58 271 62 274
rect 58 267 82 271
rect 32 259 43 263
rect 39 253 43 259
rect 78 263 82 267
rect 58 262 74 263
rect 58 260 70 262
rect 72 260 74 262
rect 58 259 74 260
rect 78 261 83 263
rect 78 259 80 261
rect 82 259 83 261
rect 58 253 62 259
rect 78 257 83 259
rect 78 255 82 257
rect 39 252 62 253
rect 39 250 41 252
rect 43 250 62 252
rect 39 249 62 250
rect 50 238 54 240
rect 50 236 51 238
rect 53 236 54 238
rect 50 231 54 236
rect 58 238 62 249
rect 66 252 82 255
rect 66 250 67 252
rect 69 251 82 252
rect 69 250 70 251
rect 66 245 70 250
rect 125 272 130 276
rect 159 275 179 276
rect 125 270 126 272
rect 128 271 151 272
rect 128 270 147 271
rect 125 269 147 270
rect 149 269 151 271
rect 125 268 151 269
rect 175 271 179 275
rect 217 279 223 285
rect 217 277 219 279
rect 221 277 223 279
rect 217 276 223 277
rect 230 276 234 278
rect 190 272 191 274
rect 175 267 187 271
rect 183 262 187 267
rect 183 260 184 262
rect 186 260 187 262
rect 66 243 67 245
rect 69 243 70 245
rect 66 241 70 243
rect 105 247 109 249
rect 105 245 106 247
rect 108 245 109 247
rect 105 240 109 245
rect 124 247 130 248
rect 124 245 126 247
rect 128 245 130 247
rect 105 238 106 240
rect 108 238 109 240
rect 58 237 91 238
rect 58 235 87 237
rect 89 235 91 237
rect 58 234 91 235
rect 50 229 51 231
rect 53 229 54 231
rect 105 229 109 238
rect 124 240 130 245
rect 183 248 187 260
rect 230 274 231 276
rect 233 274 234 276
rect 204 271 208 273
rect 204 269 205 271
rect 207 269 208 271
rect 204 263 208 269
rect 230 271 234 274
rect 230 267 254 271
rect 204 259 215 263
rect 170 245 187 248
rect 170 243 171 245
rect 173 244 187 245
rect 173 243 174 244
rect 124 238 126 240
rect 128 238 130 240
rect 124 229 130 238
rect 145 240 149 242
rect 145 238 146 240
rect 148 238 149 240
rect 145 229 149 238
rect 159 238 165 239
rect 159 236 161 238
rect 163 236 165 238
rect 159 229 165 236
rect 170 238 174 243
rect 170 236 171 238
rect 173 236 174 238
rect 170 234 174 236
rect 179 240 185 241
rect 179 238 181 240
rect 183 238 185 240
rect 179 229 185 238
rect 211 253 215 259
rect 250 263 254 267
rect 230 262 246 263
rect 230 260 242 262
rect 244 260 246 262
rect 230 259 246 260
rect 250 261 255 263
rect 250 259 252 261
rect 254 259 255 261
rect 230 253 234 259
rect 250 257 255 259
rect 250 255 254 257
rect 211 252 234 253
rect 211 250 213 252
rect 215 250 234 252
rect 211 249 234 250
rect 222 238 226 240
rect 222 236 223 238
rect 225 236 226 238
rect 222 231 226 236
rect 230 238 234 249
rect 238 252 254 255
rect 238 250 239 252
rect 241 251 254 252
rect 241 250 242 251
rect 238 245 242 250
rect 238 243 239 245
rect 241 243 242 245
rect 238 241 242 243
rect 286 274 290 285
rect 275 267 276 273
rect 286 272 287 274
rect 289 272 290 274
rect 286 270 290 272
rect 508 279 514 285
rect 466 278 486 279
rect 466 276 482 278
rect 484 276 486 278
rect 508 277 510 279
rect 512 277 514 279
rect 508 276 514 277
rect 521 276 525 278
rect 466 275 486 276
rect 275 248 276 255
rect 454 272 455 274
rect 466 271 470 275
rect 521 274 522 276
rect 524 274 525 276
rect 458 267 470 271
rect 458 262 462 267
rect 458 260 459 262
rect 461 260 462 262
rect 458 248 462 260
rect 495 271 499 273
rect 495 269 496 271
rect 498 269 499 271
rect 495 263 499 269
rect 521 271 525 274
rect 521 267 545 271
rect 495 259 506 263
rect 458 245 475 248
rect 458 244 472 245
rect 471 243 472 244
rect 474 243 475 245
rect 460 240 466 241
rect 282 238 288 239
rect 230 237 263 238
rect 230 235 259 237
rect 261 235 263 237
rect 230 234 263 235
rect 282 236 284 238
rect 286 236 288 238
rect 222 229 223 231
rect 225 229 226 231
rect 282 229 288 236
rect 460 238 462 240
rect 464 238 466 240
rect 460 229 466 238
rect 471 238 475 243
rect 502 253 506 259
rect 541 263 545 267
rect 521 262 537 263
rect 521 260 533 262
rect 535 260 537 262
rect 521 259 537 260
rect 541 261 546 263
rect 541 259 543 261
rect 545 259 546 261
rect 521 253 525 259
rect 541 257 546 259
rect 541 255 545 257
rect 502 252 525 253
rect 502 250 504 252
rect 506 250 525 252
rect 502 249 525 250
rect 471 236 472 238
rect 474 236 475 238
rect 471 234 475 236
rect 480 238 486 239
rect 480 236 482 238
rect 484 236 486 238
rect 480 229 486 236
rect 513 238 517 240
rect 513 236 514 238
rect 516 236 517 238
rect 513 231 517 236
rect 521 238 525 249
rect 529 252 545 255
rect 529 250 530 252
rect 532 251 545 252
rect 532 250 533 251
rect 529 245 533 250
rect 574 278 594 279
rect 574 276 576 278
rect 578 276 594 278
rect 574 275 594 276
rect 590 271 594 275
rect 605 272 606 274
rect 590 267 602 271
rect 598 262 602 267
rect 598 260 599 262
rect 601 260 602 262
rect 529 243 530 245
rect 532 243 533 245
rect 529 241 533 243
rect 598 248 602 260
rect 619 274 623 285
rect 619 272 620 274
rect 622 272 623 274
rect 619 270 623 272
rect 633 267 634 273
rect 647 276 651 285
rect 647 274 648 276
rect 650 274 651 276
rect 647 272 651 274
rect 585 245 602 248
rect 585 243 586 245
rect 588 244 602 245
rect 633 248 634 255
rect 588 243 589 244
rect 574 238 580 239
rect 521 237 554 238
rect 521 235 550 237
rect 552 235 554 237
rect 521 234 554 235
rect 574 236 576 238
rect 578 236 580 238
rect 513 229 514 231
rect 516 229 517 231
rect 574 229 580 236
rect 585 238 589 243
rect 585 236 586 238
rect 588 236 589 238
rect 585 234 589 236
rect 594 240 600 241
rect 594 238 596 240
rect 598 238 600 240
rect 594 229 600 238
rect 621 238 627 239
rect 621 236 623 238
rect 625 236 627 238
rect 621 229 627 236
rect 647 238 651 240
rect 647 236 648 238
rect 650 236 651 238
rect 647 231 651 236
rect 647 229 648 231
rect 650 229 651 231
rect 31 211 33 213
rect 35 211 37 213
rect 31 206 37 211
rect 31 204 33 206
rect 35 204 37 206
rect 31 203 37 204
rect 65 211 67 213
rect 69 211 71 213
rect 65 206 71 211
rect 65 204 67 206
rect 69 204 71 206
rect 65 203 71 204
rect 84 206 90 213
rect 84 204 86 206
rect 88 204 90 206
rect 84 203 90 204
rect 121 204 127 213
rect 121 202 123 204
rect 125 202 127 204
rect 121 201 127 202
rect 132 206 136 208
rect 132 204 133 206
rect 135 204 136 206
rect 132 199 136 204
rect 141 206 147 213
rect 141 204 143 206
rect 145 204 147 206
rect 141 203 147 204
rect 155 211 157 213
rect 159 211 161 213
rect 155 206 161 211
rect 155 204 157 206
rect 159 204 161 206
rect 155 203 161 204
rect 189 211 191 213
rect 193 211 195 213
rect 189 206 195 211
rect 189 204 191 206
rect 193 204 195 206
rect 189 203 195 204
rect 132 198 133 199
rect 96 187 97 194
rect 53 166 59 167
rect 53 164 55 166
rect 57 164 59 166
rect 33 159 39 160
rect 33 157 35 159
rect 37 157 39 159
rect 53 159 59 164
rect 82 170 86 172
rect 82 168 83 170
rect 85 168 86 170
rect 96 169 97 175
rect 53 157 55 159
rect 57 157 59 159
rect 82 157 86 168
rect 119 197 133 198
rect 135 197 136 199
rect 119 194 136 197
rect 119 182 123 194
rect 456 205 462 213
rect 508 211 510 213
rect 512 211 514 213
rect 456 203 458 205
rect 460 203 462 205
rect 456 202 462 203
rect 467 205 494 207
rect 467 203 468 205
rect 470 204 494 205
rect 470 203 490 204
rect 467 198 471 203
rect 488 202 490 203
rect 492 202 494 204
rect 508 206 514 211
rect 556 211 558 213
rect 560 211 562 213
rect 508 204 510 206
rect 512 204 514 206
rect 508 203 514 204
rect 533 206 537 208
rect 533 204 534 206
rect 536 204 537 206
rect 462 196 468 198
rect 470 196 471 198
rect 119 180 120 182
rect 122 180 123 182
rect 119 175 123 180
rect 119 171 131 175
rect 115 168 116 170
rect 127 167 131 171
rect 127 166 147 167
rect 127 164 143 166
rect 145 164 147 166
rect 127 163 147 164
rect 177 166 183 167
rect 177 164 179 166
rect 181 164 183 166
rect 157 159 163 160
rect 157 157 159 159
rect 161 157 163 159
rect 177 159 183 164
rect 450 189 451 195
rect 462 194 471 196
rect 462 191 466 194
rect 488 197 494 202
rect 533 199 537 204
rect 556 206 562 211
rect 556 204 558 206
rect 560 204 562 206
rect 556 203 562 204
rect 580 211 582 213
rect 584 211 586 213
rect 580 206 586 211
rect 600 211 602 213
rect 604 211 606 213
rect 580 204 582 206
rect 584 204 586 206
rect 580 203 586 204
rect 591 206 595 208
rect 591 204 592 206
rect 594 204 595 206
rect 591 200 595 204
rect 600 206 606 211
rect 651 211 652 213
rect 654 211 655 213
rect 600 204 602 206
rect 604 204 606 206
rect 614 207 647 208
rect 614 205 616 207
rect 618 205 647 207
rect 614 204 647 205
rect 600 203 606 204
rect 591 199 594 200
rect 488 195 490 197
rect 492 195 494 197
rect 488 194 494 195
rect 591 197 592 199
rect 591 195 594 197
rect 454 187 466 191
rect 454 182 458 187
rect 473 186 479 187
rect 454 180 455 182
rect 457 180 458 182
rect 454 174 458 180
rect 450 168 451 174
rect 454 170 463 174
rect 459 166 463 170
rect 582 182 583 186
rect 459 165 489 166
rect 459 163 485 165
rect 487 163 489 165
rect 459 162 489 163
rect 579 166 583 168
rect 579 164 580 166
rect 582 164 583 166
rect 177 157 179 159
rect 181 157 183 159
rect 579 159 583 164
rect 635 199 639 201
rect 635 197 636 199
rect 638 197 639 199
rect 635 192 639 197
rect 635 191 636 192
rect 623 190 636 191
rect 638 190 639 192
rect 623 187 639 190
rect 643 193 647 204
rect 651 206 655 211
rect 651 204 652 206
rect 654 204 655 206
rect 651 202 655 204
rect 643 192 666 193
rect 643 190 662 192
rect 664 190 666 192
rect 643 189 666 190
rect 623 185 627 187
rect 622 183 627 185
rect 643 183 647 189
rect 622 181 623 183
rect 625 181 627 183
rect 622 179 627 181
rect 631 182 647 183
rect 631 180 633 182
rect 635 180 647 182
rect 631 179 647 180
rect 623 175 627 179
rect 662 183 666 189
rect 662 179 673 183
rect 623 171 647 175
rect 643 168 647 171
rect 669 173 673 179
rect 669 171 670 173
rect 672 171 673 173
rect 669 169 673 171
rect 643 166 644 168
rect 646 166 647 168
rect 643 164 647 166
rect 654 165 660 166
rect 654 163 656 165
rect 658 163 660 165
rect 579 157 580 159
rect 582 157 583 159
rect 654 157 660 163
rect 45 135 51 141
rect 122 139 123 141
rect 125 139 126 141
rect 45 133 47 135
rect 49 133 51 135
rect 45 132 51 133
rect 58 132 62 134
rect 58 130 59 132
rect 61 130 62 132
rect 32 127 36 129
rect 32 125 33 127
rect 35 125 36 127
rect 32 119 36 125
rect 58 127 62 130
rect 58 123 82 127
rect 32 115 43 119
rect 39 109 43 115
rect 78 119 82 123
rect 58 118 74 119
rect 58 116 70 118
rect 72 116 74 118
rect 58 115 74 116
rect 78 117 83 119
rect 78 115 80 117
rect 82 115 83 117
rect 58 109 62 115
rect 78 113 83 115
rect 78 111 82 113
rect 39 108 62 109
rect 39 106 41 108
rect 43 106 62 108
rect 39 105 62 106
rect 50 94 54 96
rect 50 92 51 94
rect 53 92 54 94
rect 50 87 54 92
rect 58 94 62 105
rect 66 108 82 111
rect 66 106 67 108
rect 69 107 82 108
rect 69 106 70 107
rect 66 101 70 106
rect 66 99 67 101
rect 69 99 70 101
rect 66 97 70 99
rect 122 134 126 139
rect 122 132 123 134
rect 125 132 126 134
rect 122 130 126 132
rect 137 134 157 135
rect 137 132 139 134
rect 141 132 157 134
rect 137 131 157 132
rect 122 112 123 116
rect 153 127 157 131
rect 168 128 169 130
rect 153 123 165 127
rect 161 118 165 123
rect 161 116 162 118
rect 164 116 165 118
rect 111 101 114 103
rect 113 99 114 101
rect 111 98 114 99
rect 161 104 165 116
rect 148 101 165 104
rect 148 99 149 101
rect 151 100 165 101
rect 151 99 152 100
rect 99 94 105 95
rect 58 93 91 94
rect 58 91 87 93
rect 89 91 91 93
rect 58 90 91 91
rect 99 92 101 94
rect 103 92 105 94
rect 50 85 51 87
rect 53 85 54 87
rect 99 87 105 92
rect 110 94 114 98
rect 110 92 111 94
rect 113 92 114 94
rect 110 90 114 92
rect 119 94 125 95
rect 119 92 121 94
rect 123 92 125 94
rect 99 85 101 87
rect 103 85 105 87
rect 119 87 125 92
rect 119 85 121 87
rect 123 85 125 87
rect 137 94 143 95
rect 137 92 139 94
rect 141 92 143 94
rect 137 85 143 92
rect 148 94 152 99
rect 200 130 204 141
rect 189 123 190 129
rect 200 128 201 130
rect 203 128 204 130
rect 200 126 204 128
rect 451 135 455 141
rect 451 133 452 135
rect 454 133 455 135
rect 451 131 455 133
rect 493 135 497 141
rect 493 133 494 135
rect 496 133 497 135
rect 493 131 497 133
rect 523 135 553 136
rect 523 133 525 135
rect 527 133 553 135
rect 523 132 553 133
rect 189 104 190 111
rect 426 103 432 104
rect 426 101 428 103
rect 430 101 432 103
rect 148 92 149 94
rect 151 92 152 94
rect 148 90 152 92
rect 157 96 163 97
rect 157 94 159 96
rect 161 94 163 96
rect 426 96 432 101
rect 157 85 163 94
rect 196 94 202 95
rect 196 92 198 94
rect 200 92 202 94
rect 196 85 202 92
rect 426 94 428 96
rect 430 94 432 96
rect 426 85 432 94
rect 549 128 553 132
rect 493 113 494 119
rect 549 124 558 128
rect 561 124 562 130
rect 574 134 594 135
rect 574 132 576 134
rect 578 132 594 134
rect 574 131 594 132
rect 554 118 558 124
rect 554 116 555 118
rect 557 116 558 118
rect 533 111 539 112
rect 554 111 558 116
rect 546 107 558 111
rect 518 103 524 104
rect 518 101 520 103
rect 522 101 524 103
rect 518 96 524 101
rect 546 104 550 107
rect 541 102 550 104
rect 561 103 562 109
rect 590 127 594 131
rect 605 128 606 130
rect 590 123 602 127
rect 598 118 602 123
rect 598 116 599 118
rect 601 116 602 118
rect 541 100 542 102
rect 544 100 550 102
rect 518 94 520 96
rect 522 95 524 96
rect 541 95 545 100
rect 598 104 602 116
rect 619 130 623 141
rect 647 139 648 141
rect 650 139 651 141
rect 619 128 620 130
rect 622 128 623 130
rect 619 126 623 128
rect 633 123 634 129
rect 647 134 651 139
rect 647 132 648 134
rect 650 132 651 134
rect 647 130 651 132
rect 585 101 602 104
rect 585 99 586 101
rect 588 100 602 101
rect 633 104 634 111
rect 650 112 651 116
rect 588 99 589 100
rect 522 94 542 95
rect 518 93 542 94
rect 544 93 545 95
rect 518 91 545 93
rect 550 95 556 96
rect 550 93 552 95
rect 554 93 556 95
rect 550 85 556 93
rect 574 94 580 95
rect 574 92 576 94
rect 578 92 580 94
rect 574 85 580 92
rect 585 94 589 99
rect 659 101 662 103
rect 659 99 660 101
rect 659 98 662 99
rect 585 92 586 94
rect 588 92 589 94
rect 585 90 589 92
rect 594 96 600 97
rect 594 94 596 96
rect 598 94 600 96
rect 594 85 600 94
rect 621 94 627 95
rect 621 92 623 94
rect 625 92 627 94
rect 621 85 627 92
rect 648 94 654 95
rect 648 92 650 94
rect 652 92 654 94
rect 648 87 654 92
rect 659 94 663 98
rect 659 92 660 94
rect 662 92 663 94
rect 659 90 663 92
rect 668 94 674 95
rect 668 92 670 94
rect 672 92 674 94
rect 648 85 650 87
rect 652 85 654 87
rect 668 87 674 92
rect 668 85 670 87
rect 672 85 674 87
rect 31 67 33 69
rect 35 67 37 69
rect 31 62 37 67
rect 31 60 33 62
rect 35 60 37 62
rect 31 59 37 60
rect 65 67 67 69
rect 69 67 71 69
rect 65 62 71 67
rect 65 60 67 62
rect 69 60 71 62
rect 65 59 71 60
rect 82 62 88 69
rect 147 67 148 69
rect 150 67 151 69
rect 82 60 84 62
rect 86 60 88 62
rect 110 63 143 64
rect 110 61 112 63
rect 114 61 143 63
rect 110 60 143 61
rect 82 59 88 60
rect 94 43 95 50
rect 53 22 59 23
rect 53 20 55 22
rect 57 20 59 22
rect 33 15 39 16
rect 33 13 35 15
rect 37 13 39 15
rect 53 15 59 20
rect 80 26 84 28
rect 80 24 81 26
rect 83 24 84 26
rect 94 25 95 31
rect 53 13 55 15
rect 57 13 59 15
rect 80 13 84 24
rect 131 55 135 57
rect 131 53 132 55
rect 134 53 135 55
rect 131 48 135 53
rect 131 47 132 48
rect 119 46 132 47
rect 134 46 135 48
rect 119 43 135 46
rect 139 49 143 60
rect 147 62 151 67
rect 147 60 148 62
rect 150 60 151 62
rect 147 58 151 60
rect 139 48 162 49
rect 139 46 158 48
rect 160 46 162 48
rect 139 45 162 46
rect 119 41 123 43
rect 118 39 123 41
rect 139 39 143 45
rect 118 37 119 39
rect 121 37 123 39
rect 118 35 123 37
rect 127 38 143 39
rect 127 36 129 38
rect 131 36 143 38
rect 127 35 143 36
rect 119 31 123 35
rect 158 39 162 45
rect 181 60 187 69
rect 181 58 183 60
rect 185 58 187 60
rect 201 68 207 69
rect 201 66 203 68
rect 205 66 207 68
rect 201 61 207 66
rect 201 59 203 61
rect 205 59 207 61
rect 379 62 385 69
rect 431 65 435 69
rect 379 60 381 62
rect 383 60 385 62
rect 379 59 385 60
rect 201 58 207 59
rect 181 53 187 58
rect 181 51 183 53
rect 185 51 187 53
rect 181 50 187 51
rect 158 35 169 39
rect 119 27 143 31
rect 139 24 143 27
rect 165 29 169 35
rect 184 36 186 43
rect 391 43 392 50
rect 165 27 166 29
rect 168 27 169 29
rect 165 25 169 27
rect 181 25 185 27
rect 377 26 381 28
rect 139 22 140 24
rect 142 22 143 24
rect 181 23 182 25
rect 184 23 185 25
rect 377 24 378 26
rect 380 24 381 26
rect 391 25 392 31
rect 431 63 432 65
rect 434 63 435 65
rect 451 65 455 69
rect 431 61 435 63
rect 441 62 445 64
rect 441 60 442 62
rect 444 60 445 62
rect 451 63 452 65
rect 454 63 455 65
rect 503 67 504 69
rect 506 67 507 69
rect 451 61 455 63
rect 466 63 499 64
rect 466 61 468 63
rect 470 61 499 63
rect 466 60 499 61
rect 441 56 445 60
rect 424 45 429 46
rect 139 20 143 22
rect 150 21 156 22
rect 150 19 152 21
rect 154 19 156 21
rect 150 13 156 19
rect 181 13 185 23
rect 202 22 208 23
rect 202 20 204 22
rect 206 20 208 22
rect 202 13 208 20
rect 377 13 381 24
rect 424 43 425 45
rect 427 43 429 45
rect 424 42 429 43
rect 487 55 491 57
rect 487 53 488 55
rect 490 53 491 55
rect 487 48 491 53
rect 487 47 488 48
rect 475 46 488 47
rect 490 46 491 48
rect 475 43 491 46
rect 495 49 499 60
rect 503 62 507 67
rect 503 60 504 62
rect 506 60 507 62
rect 503 58 507 60
rect 534 62 540 69
rect 534 60 536 62
rect 538 60 540 62
rect 534 59 540 60
rect 545 62 549 64
rect 545 60 546 62
rect 548 60 549 62
rect 495 48 518 49
rect 495 46 514 48
rect 516 46 518 48
rect 495 45 518 46
rect 475 41 479 43
rect 474 39 479 41
rect 495 39 499 45
rect 474 37 475 39
rect 477 37 479 39
rect 474 35 479 37
rect 483 38 499 39
rect 483 36 485 38
rect 487 36 499 38
rect 483 35 499 36
rect 475 31 479 35
rect 514 39 518 45
rect 545 55 549 60
rect 554 60 560 69
rect 554 58 556 60
rect 558 58 560 60
rect 579 67 580 69
rect 582 67 583 69
rect 579 62 583 67
rect 651 67 652 69
rect 654 67 655 69
rect 614 63 647 64
rect 579 60 580 62
rect 582 60 583 62
rect 579 58 583 60
rect 614 61 616 63
rect 618 61 647 63
rect 614 60 647 61
rect 554 57 560 58
rect 545 53 546 55
rect 548 54 549 55
rect 548 53 562 54
rect 545 50 562 53
rect 514 35 525 39
rect 475 27 499 31
rect 495 24 499 27
rect 521 29 525 35
rect 521 27 522 29
rect 524 27 525 29
rect 521 25 525 27
rect 558 38 562 50
rect 558 36 559 38
rect 561 36 562 38
rect 558 31 562 36
rect 550 27 562 31
rect 495 22 496 24
rect 498 22 499 24
rect 550 23 554 27
rect 565 24 566 26
rect 534 22 554 23
rect 495 20 499 22
rect 506 21 512 22
rect 506 19 508 21
rect 510 19 512 21
rect 534 20 536 22
rect 538 20 554 22
rect 534 19 554 20
rect 506 13 512 19
rect 579 24 583 26
rect 579 22 580 24
rect 582 22 583 24
rect 579 13 583 22
rect 635 55 639 57
rect 635 53 636 55
rect 638 53 639 55
rect 635 48 639 53
rect 635 47 636 48
rect 623 46 636 47
rect 638 46 639 48
rect 623 43 639 46
rect 643 49 647 60
rect 651 62 655 67
rect 651 60 652 62
rect 654 60 655 62
rect 651 58 655 60
rect 643 48 666 49
rect 643 46 662 48
rect 664 46 666 48
rect 643 45 666 46
rect 623 41 627 43
rect 622 39 627 41
rect 643 39 647 45
rect 622 37 623 39
rect 625 37 627 39
rect 622 35 627 37
rect 631 38 647 39
rect 631 36 633 38
rect 635 36 647 38
rect 631 35 647 36
rect 623 31 627 35
rect 662 39 666 45
rect 662 35 673 39
rect 623 27 647 31
rect 643 24 647 27
rect 669 29 673 35
rect 669 27 670 29
rect 672 27 673 29
rect 669 25 673 27
rect 643 22 644 24
rect 646 22 647 24
rect 643 20 647 22
rect 654 21 660 22
rect 654 19 656 21
rect 658 19 660 21
rect 654 13 660 19
<< via1 >>
rect 40 700 42 702
rect 88 701 90 703
rect 84 676 86 678
rect 144 707 146 709
rect 116 701 118 703
rect 116 684 118 686
rect 161 698 163 700
rect 188 701 190 703
rect 105 671 107 673
rect 168 675 170 677
rect 186 667 188 669
rect 250 709 252 711
rect 274 701 276 703
rect 258 695 260 697
rect 290 698 292 700
rect 290 683 292 685
rect 325 693 327 695
rect 318 675 320 677
rect 522 684 524 686
rect 505 676 507 678
rect 552 691 554 693
rect 536 667 538 669
rect 615 701 617 703
rect 661 708 663 710
rect 661 700 663 702
rect 638 683 640 685
rect 671 684 673 686
rect 613 677 615 679
rect 96 626 98 628
rect 56 621 58 623
rect 32 605 34 607
rect 48 603 50 605
rect 84 613 86 615
rect 68 595 70 597
rect 119 620 121 622
rect 149 628 151 630
rect 120 606 122 608
rect 208 636 210 638
rect 172 620 174 622
rect 216 628 218 630
rect 164 603 166 605
rect 181 603 183 605
rect 513 628 515 630
rect 224 620 226 622
rect 505 611 507 613
rect 249 604 251 606
rect 272 605 274 607
rect 565 629 567 631
rect 533 618 535 620
rect 586 621 588 623
rect 558 603 560 605
rect 595 604 597 606
rect 603 595 605 597
rect 622 629 624 631
rect 615 604 617 606
rect 663 603 665 605
rect 40 556 42 558
rect 88 555 90 557
rect 155 564 157 566
rect 112 555 114 557
rect 147 556 149 558
rect 119 539 121 541
rect 188 540 190 542
rect 256 564 258 566
rect 224 556 226 558
rect 241 548 243 550
rect 100 531 102 533
rect 196 532 198 534
rect 223 532 225 534
rect 443 565 445 567
rect 537 556 539 558
rect 459 549 461 551
rect 487 548 489 550
rect 567 556 569 558
rect 559 540 561 542
rect 529 534 531 536
rect 646 556 648 558
rect 619 548 621 550
rect 605 536 607 538
rect 638 539 640 541
rect 594 532 596 534
rect 655 535 657 537
rect 56 477 58 479
rect 56 469 58 471
rect 32 459 34 461
rect 128 484 130 486
rect 29 451 31 453
rect 76 459 78 461
rect 96 460 98 462
rect 68 451 70 453
rect 136 451 138 453
rect 200 492 202 494
rect 220 485 222 487
rect 191 460 193 462
rect 251 481 253 483
rect 228 459 230 461
rect 498 493 500 495
rect 543 484 545 486
rect 489 460 491 462
rect 511 460 513 462
rect 620 484 622 486
rect 575 476 577 478
rect 536 468 538 470
rect 558 468 560 470
rect 603 469 605 471
rect 663 460 665 462
rect 615 452 617 454
rect 29 413 31 415
rect 57 413 59 415
rect 48 400 50 402
rect 92 413 94 415
rect 91 396 93 398
rect 68 382 70 384
rect 141 410 143 412
rect 117 391 119 393
rect 180 404 182 406
rect 149 387 151 389
rect 202 399 204 401
rect 170 388 172 390
rect 216 410 218 412
rect 232 403 234 405
rect 268 413 270 415
rect 244 391 246 393
rect 276 396 278 398
rect 329 413 331 415
rect 312 404 314 406
rect 435 404 437 406
rect 289 380 291 382
rect 321 388 323 390
rect 450 413 452 415
rect 418 387 420 389
rect 471 413 473 415
rect 498 413 500 415
rect 491 395 493 397
rect 471 387 473 389
rect 523 390 525 392
rect 540 390 542 392
rect 554 404 556 406
rect 586 408 588 410
rect 635 421 637 423
rect 612 404 614 406
rect 571 387 573 389
rect 595 389 597 391
rect 655 412 657 414
rect 639 387 641 389
rect 650 384 652 386
rect 53 344 55 346
rect 64 341 66 343
rect 48 316 50 318
rect 108 339 110 341
rect 132 341 134 343
rect 91 324 93 326
rect 68 307 70 309
rect 117 320 119 322
rect 149 324 151 326
rect 163 338 165 340
rect 76 307 78 309
rect 180 338 182 340
rect 232 341 234 343
rect 212 333 214 335
rect 205 315 207 317
rect 232 315 234 317
rect 285 341 287 343
rect 253 315 255 317
rect 382 340 384 342
rect 414 348 416 350
rect 268 324 270 326
rect 391 324 393 326
rect 374 315 376 317
rect 427 332 429 334
rect 459 337 461 339
rect 435 315 437 317
rect 471 325 473 327
rect 487 318 489 320
rect 533 340 535 342
rect 501 329 503 331
rect 554 341 556 343
rect 523 324 525 326
rect 586 337 588 339
rect 562 318 564 320
rect 635 346 637 348
rect 612 332 614 334
rect 611 315 613 317
rect 655 328 657 330
rect 646 315 648 317
rect 674 315 676 317
rect 88 276 90 278
rect 40 268 42 270
rect 100 259 102 261
rect 145 260 147 262
rect 167 260 169 262
rect 128 252 130 254
rect 83 244 85 246
rect 192 268 194 270
rect 214 268 216 270
rect 160 244 162 246
rect 205 235 207 237
rect 280 268 282 270
rect 475 269 477 271
rect 280 244 282 246
rect 452 247 454 249
rect 512 268 514 270
rect 483 243 485 245
rect 503 236 505 238
rect 567 277 569 279
rect 635 277 637 279
rect 607 268 609 270
rect 627 269 629 271
rect 674 277 676 279
rect 575 244 577 246
rect 671 269 673 271
rect 647 259 649 261
rect 647 251 649 253
rect 48 193 50 195
rect 109 196 111 198
rect 65 189 67 191
rect 98 192 100 194
rect 84 180 86 182
rect 57 172 59 174
rect 174 194 176 196
rect 144 188 146 190
rect 136 172 138 174
rect 216 180 218 182
rect 166 172 168 174
rect 480 196 482 198
rect 507 196 509 198
rect 603 197 605 199
rect 462 180 464 182
rect 479 172 481 174
rect 447 164 449 166
rect 515 188 517 190
rect 584 189 586 191
rect 556 172 558 174
rect 591 173 593 175
rect 548 164 550 166
rect 615 173 617 175
rect 663 172 665 174
rect 40 125 42 127
rect 88 124 90 126
rect 81 99 83 101
rect 100 133 102 135
rect 108 124 110 126
rect 145 125 147 127
rect 117 107 119 109
rect 170 110 172 112
rect 138 99 140 101
rect 431 123 433 125
rect 454 124 456 126
rect 198 117 200 119
rect 479 108 481 110
rect 190 100 192 102
rect 522 125 524 127
rect 539 125 541 127
rect 487 100 489 102
rect 531 108 533 110
rect 495 92 497 94
rect 583 122 585 124
rect 554 100 556 102
rect 584 108 586 110
rect 635 133 637 135
rect 619 115 621 117
rect 655 125 657 127
rect 671 123 673 125
rect 647 107 649 109
rect 607 102 609 104
rect 90 51 92 53
rect 32 44 34 46
rect 65 45 67 47
rect 42 28 44 30
rect 42 20 44 22
rect 88 27 90 29
rect 167 61 169 63
rect 151 37 153 39
rect 198 52 200 54
rect 190 44 192 46
rect 385 53 387 55
rect 378 35 380 37
rect 413 45 415 47
rect 413 30 415 32
rect 445 33 447 35
rect 429 27 431 29
rect 453 19 455 21
rect 517 61 519 63
rect 535 53 537 55
rect 598 57 600 59
rect 515 27 517 29
rect 542 30 544 32
rect 587 44 589 46
rect 587 27 589 29
rect 559 21 561 23
rect 619 52 621 54
rect 615 27 617 29
rect 663 28 665 30
<< via2 >>
rect 266 701 268 703
rect 32 590 34 592
rect 299 698 301 700
rect 161 694 163 696
rect 32 463 34 465
rect 96 642 98 644
rect 115 620 117 622
rect 125 606 127 608
rect 153 642 155 644
rect 288 642 290 644
rect 164 582 166 584
rect 181 606 183 608
rect 296 597 298 599
rect 288 589 290 591
rect 172 582 174 584
rect 108 572 110 574
rect 85 563 87 565
rect 321 548 323 550
rect 100 498 102 500
rect 223 528 225 530
rect 100 484 102 486
rect 223 485 225 487
rect 260 485 262 487
rect 56 459 58 461
rect 72 459 74 461
rect 221 459 223 461
rect 72 436 74 438
rect 296 436 298 438
rect 100 426 102 428
rect 276 426 278 428
rect 108 418 110 420
rect 64 374 66 376
rect 68 332 70 334
rect 48 312 50 314
rect 132 418 134 420
rect 172 410 174 412
rect 206 410 208 412
rect 155 387 157 389
rect 132 374 134 376
rect 149 354 151 356
rect 221 374 223 376
rect 232 354 234 356
rect 227 333 229 335
rect 76 282 78 284
rect 214 282 216 284
rect 136 158 138 160
rect 227 218 229 220
rect 198 158 200 160
rect 208 142 210 144
rect 136 133 138 135
rect 32 86 34 88
rect 198 112 200 114
rect 321 167 323 169
rect 329 158 331 160
rect 374 570 376 572
rect 382 561 384 563
rect 487 642 489 644
rect 505 616 507 618
rect 671 642 673 644
rect 567 595 569 597
rect 495 586 497 588
rect 505 570 507 572
rect 476 510 478 512
rect 567 570 569 572
rect 476 395 478 397
rect 471 374 473 376
rect 482 354 484 356
rect 554 374 556 376
rect 571 354 573 356
rect 548 341 550 343
rect 497 318 499 320
rect 531 318 533 320
rect 571 310 573 312
rect 655 416 657 418
rect 635 396 637 398
rect 639 354 641 356
rect 595 310 597 312
rect 427 302 429 304
rect 603 302 605 304
rect 407 292 409 294
rect 631 292 633 294
rect 482 269 484 271
rect 631 269 633 271
rect 647 269 649 271
rect 443 243 445 245
rect 480 243 482 245
rect 603 244 605 246
rect 480 200 482 202
rect 603 230 605 232
rect 382 180 384 182
rect 216 86 218 88
rect 618 165 620 167
rect 595 156 597 158
rect 531 146 533 148
rect 415 139 417 141
rect 407 131 409 133
rect 522 122 524 124
rect 539 146 541 148
rect 415 86 417 88
rect 550 86 552 88
rect 578 122 580 124
rect 588 108 590 110
rect 607 86 609 88
rect 671 265 673 267
rect 542 34 544 36
rect 404 30 406 32
rect 671 138 673 140
rect 437 27 439 29
<< labels >>
rlabel space 24 0 214 149 1 PART1
rlabel space 24 149 270 298 1 PART2
rlabel space 24 298 346 437 1 PART5
rlabel space 24 437 259 581 1 PART3
rlabel space 27 581 283 725 1 PART4
rlabel alu1 182 43 182 43 1 add_sub
rlabel alu1 122 109 122 109 1 A0
rlabel alu1 112 32 112 32 1 S0
rlabel alu1 33 95 33 95 1 B0
rlabel alu1 33 238 33 238 1 B1
rlabel alu1 101 270 101 270 1 A1
rlabel alu1 261 266 261 266 1 S1
rlabel alu1 34 525 34 525 1 B2
rlabel alu1 124 540 124 540 1 A2
rlabel alu1 153 467 153 467 1 S2
rlabel alu1 34 671 34 671 1 B3
rlabel alu1 114 688 114 688 1 A3
rlabel alu1 237 698 237 698 1 S3
rlabel alu1 108 9 108 9 1 Vss
rlabel alu1 105 76 105 76 1 Vdd
rlabel alu1 100 150 100 150 1 Vss
rlabel alu1 101 222 101 222 1 Vdd
rlabel alu1 100 293 100 293 1 Vss
rlabel alu1 105 365 105 365 1 Vdd
rlabel alu1 105 433 105 433 1 Vss
rlabel alu1 105 509 105 509 1 Vdd
rlabel alu1 101 580 101 580 1 Vss
rlabel alu1 101 654 101 654 1 Vdd
rlabel alu1 96 721 96 721 1 Vss
rlabel alu1 77 329 77 329 1 co1
rlabel alu1 281 289 281 289 8 vss
rlabel alu1 281 225 281 225 8 vdd
rlabel space 24 77 99 149 1 xor2v0x1
rlabel space 24 0 75 77 1 nr2v0x2
rlabel space 75 0 102 77 1 iv1v0x1
rlabel space 131 77 179 149 1 an2v0x1
rlabel space 99 77 131 149 1 nd2v0x2
rlabel space 102 0 179 77 1 xor2v0x1
rlabel space 180 77 211 147 1 iv1v0x1
rlabel space 180 5 211 73 1 iv1v0x3
rlabel space 491 581 681 730 5 PART1
rlabel space 435 432 681 581 5 PART2
rlabel space 359 293 681 432 5 PART5
rlabel space 446 149 681 293 5 PART3
rlabel space 422 5 678 149 5 PART4
rlabel alu1 597 721 597 721 5 Vss
rlabel alu1 600 654 600 654 5 Vdd
rlabel alu1 605 580 605 580 5 Vss
rlabel alu1 604 508 604 508 5 Vdd
rlabel alu1 605 437 605 437 5 Vss
rlabel alu1 600 365 600 365 5 Vdd
rlabel alu1 600 297 600 297 5 Vss
rlabel alu1 600 221 600 221 5 Vdd
rlabel alu1 604 150 604 150 5 Vss
rlabel alu1 604 76 604 76 5 Vdd
rlabel alu1 609 9 609 9 5 Vss
rlabel alu1 593 698 593 698 5 S4
rlabel alu1 583 621 583 621 5 A4
rlabel alu1 672 635 672 635 5 B4
rlabel alu1 604 460 604 460 5 A5
rlabel alu1 672 492 672 492 5 B5
rlabel alu1 444 464 444 464 5 S5
rlabel alu1 628 401 628 401 5 Cout
rlabel alu1 552 263 552 263 5 S6
rlabel alu1 671 205 671 205 5 B6
rlabel alu1 581 190 581 190 5 A6
rlabel alu1 591 42 591 42 5 A7
rlabel alu1 671 59 671 59 5 B7
rlabel alu1 468 32 468 32 5 S7
rlabel alu1 452 577 452 577 8 vss
rlabel alu1 452 513 452 513 8 vdd
rlabel space 27 223 95 294 1 xor2v0x1
rlabel space 96 223 155 294 1 nd2v0x3
rlabel space 27 151 80 220 1 nr2v0x2
rlabel space 81 152 107 220 1 iv1v0x1
rlabel space 156 223 202 294 1 an2v0x1
rlabel space 203 223 266 294 1 xor2v0x1
rlabel space 108 152 151 220 1 an2v0x1
rlabel space 152 152 203 220 1 nr2v0x2
rlabel space 15 85 15 85 3 SUM0
rlabel space 12 225 12 225 3 SUM1
rlabel space 0 365 0 365 3 CARRY_FORWARD
rlabel space 167 369 211 430 1 an2v0x1
rlabel space 115 369 161 430 1 an2v0x1
rlabel space 62 369 105 430 1 an2v0x1
rlabel space 212 369 238 430 1 iv1v0x1
rlabel space 239 369 282 430 1 an2v0x1
rlabel ab 285 369 336 430 1 an3v0x1
rlabel ab 74 300 125 359 1 an3v0x1
rlabel space 127 300 170 359 1 an2v0x1
rlabel space 177 300 220 359 1 an2v0x1
rlabel space 246 300 289 359 1 an2v0x1
rlabel ab 221 300 244 359 1 iv1v0x1
rlabel space 27 300 72 359 1 nd3v0x1
rlabel space 28 369 60 430 1 nd2v0x1
rlabel space 62 442 89 505 1 iv1v0x1
rlabel space 93 442 138 505 1 an2v0x1
rlabel ab 217 441 257 504 1 an2v0x1
rlabel space 141 442 213 505 1 xor2v0x1
rlabel space 29 509 95 576 1 xor2v0x1
rlabel space 97 514 131 576 1 nd2v0x2
rlabel space 139 514 206 576 1 nr3v0x1
rlabel space 28 441 61 505 1 nr2v0x1
rlabel ab 271 227 290 293 1 iv1v0x1
rlabel ab 210 515 259 578 1 an3v0x1
rlabel space 64 591 90 647 1 iv1v0x1
rlabel space 131 656 174 722 1 an2v0x1
rlabel ab 93 591 132 647 1 an2v0x1
rlabel space 305 656 333 723 1 iv1v0x1
rlabel ab 29 656 92 722 1 xor2v0x1
rlabel space 177 656 245 722 1 xor2v0x1
rlabel ab 203 586 281 651 1 nr4v0x1
rlabel ab 98 656 128 722 1 nr2v0x1
rlabel ab 29 586 61 648 1 nd2v0x2
rlabel ab 137 591 195 646 1 an3v0x1
rlabel ab 247 656 302 722 1 nd4v0x1
rlabel space 12 465 12 465 1 SUM2
rlabel space 8 657 8 657 1 SUM3
<< end >>
