magic
tech scmos
timestamp 1554063197
<< ab >>
rect 78 1116 142 1188
rect 146 1116 178 1188
rect 182 1116 222 1188
rect 226 1116 292 1188
rect 296 1116 352 1188
rect 356 1116 380 1188
rect 560 1156 563 1193
rect 560 1117 563 1155
rect 564 1152 596 1188
rect 564 1148 598 1152
rect 564 1117 596 1148
rect 565 1116 597 1117
rect 602 1116 666 1188
rect 673 1116 745 1188
rect 78 1044 110 1116
rect 114 1056 138 1116
rect 142 1056 182 1116
rect 186 1056 334 1116
rect 563 1108 565 1116
rect 112 1052 334 1056
rect 114 1044 138 1052
rect 142 1044 182 1052
rect 186 1044 334 1052
rect 567 1044 591 1116
rect 599 1044 639 1116
rect 645 1044 677 1116
rect 681 1044 745 1116
rect 78 1005 142 1044
rect 146 1005 178 1044
rect 78 1001 178 1005
rect 78 972 144 1001
rect 146 972 178 1001
rect 182 972 184 1044
rect 186 1006 250 1044
rect 254 1006 308 1044
rect 186 1002 308 1006
rect 186 972 250 1002
rect 254 972 308 1002
rect 509 972 533 1044
rect 535 1036 572 1044
rect 535 972 572 980
rect 573 972 621 1044
rect 625 972 665 1044
rect 669 1041 693 1044
rect 669 973 670 1041
rect 671 973 694 1041
rect 669 972 693 973
rect 697 972 745 1044
rect 78 917 110 972
rect 77 913 110 917
rect 78 899 110 913
rect 114 900 138 972
rect 140 939 182 972
rect 142 902 182 939
rect 142 900 184 902
rect 198 900 262 972
rect 266 902 306 972
rect 266 900 308 902
rect 509 900 573 972
rect 577 900 617 972
rect 621 900 677 972
rect 681 900 745 972
rect 79 879 111 899
rect 77 873 111 879
rect 79 829 111 873
rect 114 829 154 900
rect 158 892 213 900
rect 163 836 203 892
rect 156 830 203 836
rect 205 830 213 836
rect 216 830 256 900
rect 260 830 261 900
rect 73 828 154 829
rect 158 828 214 830
rect 218 828 258 830
rect 262 828 286 900
rect 290 828 330 900
rect 334 828 390 900
rect 485 899 509 900
rect 513 899 553 900
rect 484 828 524 899
rect 529 861 553 899
rect 529 828 554 861
rect 557 828 597 900
rect 601 898 641 900
rect 645 898 701 900
rect 599 828 601 898
rect 605 828 645 898
rect 647 831 701 898
rect 705 831 745 900
rect 647 828 750 831
rect 73 825 176 828
rect 78 756 118 825
rect 122 758 176 825
rect 178 758 218 828
rect 222 758 224 828
rect 122 756 178 758
rect 182 756 222 758
rect 226 756 266 828
rect 269 795 294 828
rect 270 757 294 795
rect 299 757 339 828
rect 270 756 310 757
rect 314 756 338 757
rect 433 756 489 828
rect 493 756 533 828
rect 537 756 561 828
rect 565 826 605 828
rect 609 826 665 828
rect 669 827 750 828
rect 562 756 563 826
rect 567 756 607 826
rect 610 820 618 826
rect 620 820 667 826
rect 620 764 660 820
rect 610 756 665 764
rect 669 756 709 827
rect 712 783 744 827
rect 712 777 746 783
rect 712 757 744 777
rect 78 684 142 756
rect 146 684 202 756
rect 206 684 246 756
rect 250 684 314 756
rect 318 684 342 756
rect 515 754 557 756
rect 517 684 557 754
rect 561 684 625 756
rect 639 754 681 756
rect 641 717 681 754
rect 641 684 683 717
rect 685 684 709 756
rect 713 743 745 757
rect 713 739 746 743
rect 713 684 745 739
rect 78 612 126 684
rect 130 683 154 684
rect 129 615 152 683
rect 153 615 154 683
rect 130 612 154 615
rect 158 612 198 684
rect 202 612 250 684
rect 515 654 569 684
rect 573 654 637 684
rect 515 650 637 654
rect 515 612 569 650
rect 573 612 637 650
rect 639 612 641 684
rect 645 655 677 684
rect 679 655 745 684
rect 645 651 745 655
rect 645 612 677 651
rect 681 612 745 651
rect 78 540 142 612
rect 146 540 178 612
rect 184 540 224 612
rect 232 540 256 612
rect 489 604 637 612
rect 641 604 681 612
rect 685 604 709 612
rect 489 600 711 604
rect 258 540 260 548
rect 489 540 637 600
rect 641 540 681 600
rect 685 540 709 600
rect 713 540 745 612
rect 78 468 150 540
rect 157 468 221 540
rect 226 539 258 540
rect 227 508 259 539
rect 225 504 259 508
rect 227 468 259 504
rect 260 501 263 539
rect 260 463 263 500
rect 443 468 467 540
rect 471 468 527 540
rect 531 468 597 540
rect 601 468 641 540
rect 645 468 677 540
rect 681 468 745 540
rect 3 285 99 365
rect 3 281 102 285
rect 3 264 99 281
rect 103 264 199 365
rect 203 265 299 365
rect 303 289 399 365
rect 403 293 499 365
rect 503 293 599 365
rect 603 293 699 365
rect 703 293 799 365
rect 405 289 501 293
rect 505 289 601 293
rect 303 285 601 289
rect 3 260 102 264
rect 103 260 202 264
rect 203 261 302 265
rect 3 5 99 260
rect 103 120 199 260
rect 103 116 202 120
rect 103 5 199 116
rect 203 5 299 261
rect 303 237 399 285
rect 405 237 501 285
rect 505 237 601 285
rect 605 265 701 293
rect 605 261 704 265
rect 605 237 701 261
rect 303 233 701 237
rect 303 5 399 233
rect 405 211 501 233
rect 505 211 601 233
rect 605 211 701 233
rect 705 211 801 293
rect 400 209 801 211
rect 405 77 501 209
rect 505 77 601 209
rect 605 77 701 209
rect 705 77 801 209
rect 806 109 820 189
rect 403 5 499 77
rect 503 5 599 77
rect 603 5 699 77
rect 703 5 799 77
rect -14 -95 82 -23
rect 92 -87 188 -23
rect 92 -95 197 -87
rect 198 -95 294 -23
rect 304 -87 400 -23
rect 295 -95 400 -87
rect 410 -95 506 -23
rect 516 -95 612 -23
rect 622 -87 718 -23
rect 728 -31 930 -23
rect 728 -87 824 -31
rect 622 -95 824 -87
rect 825 -95 833 -87
rect 834 -95 930 -31
<< nwell >>
rect 73 1116 385 1156
rect 73 1076 336 1116
rect 560 1076 750 1156
rect 73 967 311 1012
rect 73 932 308 967
rect 504 932 750 1012
rect 73 823 390 868
rect 480 833 750 868
rect 73 788 343 823
rect 428 788 750 833
rect 73 679 347 724
rect 515 689 750 724
rect 73 644 255 679
rect 512 644 750 689
rect 73 500 263 580
rect 487 540 750 580
rect 438 500 750 540
rect -2 298 804 333
rect -2 253 820 298
rect -2 109 820 189
rect -2 0 804 45
rect -19 -63 935 -18
<< pwell >>
rect 73 1188 379 1193
rect 73 1156 385 1188
rect 560 1156 750 1193
rect 73 1044 336 1076
rect 560 1049 750 1076
rect 73 1039 335 1044
rect 73 1012 311 1039
rect 504 1012 750 1049
rect 73 905 308 932
rect 504 905 750 932
rect 73 868 390 905
rect 480 868 750 905
rect 73 761 343 788
rect 73 724 347 761
rect 428 751 750 788
rect 515 724 750 751
rect 73 617 255 644
rect 512 617 750 644
rect 73 580 263 617
rect 488 612 750 617
rect 487 580 750 612
rect 73 463 263 500
rect 438 468 750 500
rect 444 463 750 468
rect -2 333 804 370
rect -2 189 820 253
rect -2 72 820 109
rect -2 45 804 72
rect -19 -100 935 -63
<< poly >>
rect 90 1184 115 1186
rect 90 1176 92 1184
rect 103 1176 105 1180
rect 113 1176 115 1184
rect 123 1179 125 1184
rect 130 1179 132 1184
rect 87 1174 92 1176
rect 87 1171 89 1174
rect 156 1176 158 1181
rect 167 1173 169 1177
rect 191 1173 193 1177
rect 204 1175 206 1180
rect 211 1175 213 1180
rect 238 1184 263 1186
rect 238 1176 240 1184
rect 251 1176 253 1180
rect 261 1176 263 1184
rect 271 1179 273 1184
rect 278 1179 280 1184
rect 311 1182 313 1186
rect 318 1182 320 1186
rect 325 1182 327 1186
rect 332 1182 334 1186
rect 103 1164 105 1167
rect 96 1162 105 1164
rect 113 1163 115 1167
rect 123 1164 125 1167
rect 87 1154 89 1162
rect 96 1160 98 1162
rect 100 1160 105 1162
rect 96 1158 105 1160
rect 121 1162 125 1164
rect 121 1159 123 1162
rect 103 1154 105 1158
rect 117 1157 123 1159
rect 130 1158 132 1167
rect 156 1159 158 1168
rect 167 1162 169 1165
rect 235 1174 240 1176
rect 235 1171 237 1174
rect 165 1160 171 1162
rect 117 1155 119 1157
rect 121 1155 123 1157
rect 84 1152 97 1154
rect 103 1152 113 1154
rect 117 1153 123 1155
rect 84 1151 86 1152
rect 80 1149 86 1151
rect 95 1149 97 1152
rect 111 1149 113 1152
rect 121 1149 123 1153
rect 127 1156 133 1158
rect 127 1154 129 1156
rect 131 1154 133 1156
rect 127 1152 133 1154
rect 155 1157 161 1159
rect 155 1155 157 1157
rect 159 1155 161 1157
rect 155 1153 161 1155
rect 165 1158 167 1160
rect 169 1158 171 1160
rect 165 1156 171 1158
rect 191 1159 193 1164
rect 204 1159 206 1164
rect 191 1157 197 1159
rect 131 1149 133 1152
rect 158 1150 160 1153
rect 165 1150 167 1156
rect 191 1155 193 1157
rect 195 1155 197 1157
rect 191 1153 197 1155
rect 201 1157 207 1159
rect 201 1155 203 1157
rect 205 1155 207 1157
rect 201 1153 207 1155
rect 80 1147 82 1149
rect 84 1147 86 1149
rect 80 1145 86 1147
rect 111 1127 113 1131
rect 121 1127 123 1131
rect 95 1118 97 1122
rect 191 1149 193 1153
rect 201 1142 203 1153
rect 211 1151 213 1164
rect 251 1164 253 1167
rect 244 1162 253 1164
rect 261 1163 263 1167
rect 271 1164 273 1167
rect 235 1154 237 1162
rect 244 1160 246 1162
rect 248 1160 253 1162
rect 244 1158 253 1160
rect 269 1162 273 1164
rect 269 1159 271 1162
rect 251 1154 253 1158
rect 265 1157 271 1159
rect 278 1158 280 1167
rect 614 1184 639 1186
rect 365 1171 367 1176
rect 574 1172 576 1177
rect 584 1172 586 1177
rect 614 1176 616 1184
rect 627 1176 629 1180
rect 637 1176 639 1184
rect 647 1179 649 1184
rect 654 1179 656 1184
rect 722 1182 724 1186
rect 732 1182 734 1186
rect 611 1174 616 1176
rect 611 1171 613 1174
rect 682 1171 684 1176
rect 627 1164 629 1167
rect 620 1162 629 1164
rect 637 1163 639 1167
rect 647 1164 649 1167
rect 311 1159 313 1162
rect 265 1155 267 1157
rect 269 1155 271 1157
rect 232 1152 245 1154
rect 251 1152 261 1154
rect 265 1153 271 1155
rect 232 1151 234 1152
rect 211 1149 217 1151
rect 211 1147 213 1149
rect 215 1147 217 1149
rect 211 1145 217 1147
rect 228 1149 234 1151
rect 243 1149 245 1152
rect 259 1149 261 1152
rect 269 1149 271 1153
rect 275 1156 281 1158
rect 275 1154 277 1156
rect 279 1154 281 1156
rect 275 1152 281 1154
rect 279 1149 281 1152
rect 305 1157 313 1159
rect 305 1155 307 1157
rect 309 1156 313 1157
rect 309 1155 311 1156
rect 305 1153 311 1155
rect 228 1147 230 1149
rect 232 1147 234 1149
rect 228 1145 234 1147
rect 211 1142 213 1145
rect 191 1127 193 1131
rect 201 1124 203 1129
rect 211 1124 213 1129
rect 131 1118 133 1122
rect 158 1118 160 1122
rect 165 1118 167 1122
rect 259 1127 261 1131
rect 269 1127 271 1131
rect 243 1118 245 1122
rect 305 1143 307 1153
rect 318 1152 320 1162
rect 325 1152 327 1162
rect 332 1159 334 1162
rect 365 1159 367 1162
rect 332 1157 343 1159
rect 335 1155 339 1157
rect 341 1155 343 1157
rect 335 1153 343 1155
rect 365 1157 371 1159
rect 365 1155 367 1157
rect 369 1155 371 1157
rect 365 1153 371 1155
rect 574 1154 576 1162
rect 584 1158 586 1162
rect 584 1156 594 1158
rect 584 1154 590 1156
rect 592 1154 594 1156
rect 611 1154 613 1162
rect 620 1160 622 1162
rect 624 1160 629 1162
rect 620 1158 629 1160
rect 645 1162 649 1164
rect 645 1159 647 1162
rect 627 1154 629 1158
rect 641 1157 647 1159
rect 654 1158 656 1167
rect 706 1165 712 1167
rect 706 1163 708 1165
rect 710 1163 712 1165
rect 682 1159 684 1162
rect 706 1161 712 1163
rect 641 1155 643 1157
rect 645 1155 647 1157
rect 315 1150 321 1152
rect 315 1148 317 1150
rect 319 1148 321 1150
rect 315 1146 321 1148
rect 325 1150 331 1152
rect 325 1148 327 1150
rect 329 1148 331 1150
rect 325 1146 331 1148
rect 315 1143 317 1146
rect 325 1143 327 1146
rect 335 1143 337 1153
rect 365 1150 367 1153
rect 574 1152 594 1154
rect 608 1152 621 1154
rect 627 1152 637 1154
rect 641 1153 647 1155
rect 574 1147 576 1152
rect 584 1147 586 1152
rect 608 1151 610 1152
rect 604 1149 610 1151
rect 619 1149 621 1152
rect 635 1149 637 1152
rect 645 1149 647 1153
rect 651 1156 657 1158
rect 651 1154 653 1156
rect 655 1154 657 1156
rect 651 1152 657 1154
rect 655 1149 657 1152
rect 682 1157 688 1159
rect 682 1155 684 1157
rect 686 1155 688 1157
rect 682 1153 688 1155
rect 682 1150 684 1153
rect 604 1147 606 1149
rect 608 1147 610 1149
rect 365 1127 367 1132
rect 279 1118 281 1122
rect 305 1121 307 1126
rect 315 1121 317 1126
rect 325 1121 327 1126
rect 335 1121 337 1126
rect 604 1145 610 1147
rect 584 1127 586 1131
rect 574 1119 576 1123
rect 635 1127 637 1131
rect 645 1127 647 1131
rect 619 1118 621 1122
rect 710 1149 712 1161
rect 722 1159 724 1167
rect 732 1164 734 1167
rect 717 1157 724 1159
rect 728 1162 734 1164
rect 728 1160 730 1162
rect 732 1161 734 1162
rect 732 1160 736 1161
rect 728 1158 736 1160
rect 717 1155 719 1157
rect 721 1155 724 1157
rect 717 1154 724 1155
rect 717 1152 729 1154
rect 717 1149 719 1152
rect 727 1149 729 1152
rect 734 1149 736 1158
rect 682 1127 684 1132
rect 655 1118 657 1122
rect 710 1118 712 1122
rect 717 1118 719 1122
rect 727 1118 729 1122
rect 734 1118 736 1122
rect 87 1110 89 1114
rect 97 1110 99 1114
rect 123 1100 125 1105
rect 151 1101 153 1105
rect 161 1103 163 1108
rect 171 1103 173 1108
rect 87 1079 89 1086
rect 97 1083 99 1086
rect 97 1081 108 1083
rect 195 1102 197 1107
rect 205 1102 207 1107
rect 215 1102 217 1107
rect 267 1108 269 1113
rect 274 1108 276 1113
rect 281 1108 283 1113
rect 288 1108 290 1113
rect 97 1079 104 1081
rect 106 1079 108 1081
rect 87 1077 93 1079
rect 87 1075 89 1077
rect 91 1075 93 1077
rect 87 1073 93 1075
rect 97 1077 108 1079
rect 123 1079 125 1082
rect 151 1079 153 1083
rect 161 1079 163 1090
rect 171 1087 173 1090
rect 171 1085 177 1087
rect 171 1083 173 1085
rect 175 1083 177 1085
rect 227 1101 229 1106
rect 171 1081 177 1083
rect 123 1077 129 1079
rect 90 1070 92 1073
rect 97 1070 99 1077
rect 123 1075 125 1077
rect 127 1075 129 1077
rect 123 1073 129 1075
rect 151 1077 157 1079
rect 151 1075 153 1077
rect 155 1075 157 1077
rect 151 1073 157 1075
rect 161 1077 167 1079
rect 161 1075 163 1077
rect 165 1075 167 1077
rect 161 1073 167 1075
rect 123 1070 125 1073
rect 151 1068 153 1073
rect 164 1068 166 1073
rect 171 1068 173 1081
rect 195 1079 197 1084
rect 205 1079 207 1089
rect 215 1086 217 1089
rect 215 1084 221 1086
rect 215 1082 217 1084
rect 219 1082 221 1084
rect 215 1080 221 1082
rect 195 1077 201 1079
rect 195 1075 197 1077
rect 199 1075 201 1077
rect 195 1073 201 1075
rect 205 1077 211 1079
rect 205 1075 207 1077
rect 209 1075 211 1077
rect 205 1073 211 1075
rect 195 1069 197 1073
rect 208 1069 210 1073
rect 215 1069 217 1080
rect 227 1079 229 1088
rect 656 1110 658 1114
rect 666 1110 668 1114
rect 690 1110 692 1114
rect 298 1101 300 1105
rect 305 1101 307 1105
rect 312 1101 314 1105
rect 319 1101 321 1105
rect 580 1100 582 1105
rect 608 1101 610 1105
rect 618 1103 620 1108
rect 628 1103 630 1108
rect 267 1080 269 1083
rect 227 1077 233 1079
rect 227 1075 229 1077
rect 231 1075 233 1077
rect 222 1073 233 1075
rect 256 1078 269 1080
rect 256 1076 258 1078
rect 260 1076 265 1078
rect 256 1074 265 1076
rect 222 1069 224 1073
rect 123 1056 125 1061
rect 151 1055 153 1059
rect 90 1046 92 1050
rect 97 1046 99 1050
rect 164 1052 166 1057
rect 171 1052 173 1057
rect 195 1055 197 1060
rect 263 1062 265 1074
rect 274 1073 276 1083
rect 281 1080 283 1083
rect 288 1080 290 1083
rect 298 1080 300 1083
rect 281 1077 284 1080
rect 288 1078 300 1080
rect 271 1071 277 1073
rect 271 1069 273 1071
rect 275 1069 277 1071
rect 271 1067 277 1069
rect 282 1071 284 1077
rect 282 1069 288 1071
rect 282 1067 284 1069
rect 286 1067 288 1069
rect 273 1062 275 1067
rect 282 1065 288 1067
rect 285 1062 287 1065
rect 295 1062 297 1078
rect 305 1071 307 1083
rect 312 1074 314 1083
rect 319 1080 321 1083
rect 319 1078 327 1080
rect 580 1079 582 1082
rect 321 1076 323 1078
rect 325 1076 327 1078
rect 321 1074 327 1076
rect 576 1077 582 1079
rect 576 1075 578 1077
rect 580 1075 582 1077
rect 301 1069 307 1071
rect 301 1067 303 1069
rect 305 1067 307 1069
rect 311 1072 317 1074
rect 576 1073 582 1075
rect 311 1070 313 1072
rect 315 1070 317 1072
rect 580 1070 582 1073
rect 608 1079 610 1083
rect 618 1079 620 1090
rect 628 1087 630 1090
rect 628 1085 634 1087
rect 628 1083 630 1085
rect 632 1083 634 1085
rect 656 1083 658 1086
rect 628 1081 634 1083
rect 647 1081 658 1083
rect 608 1077 614 1079
rect 608 1075 610 1077
rect 612 1075 614 1077
rect 608 1073 614 1075
rect 618 1077 624 1079
rect 618 1075 620 1077
rect 622 1075 624 1077
rect 618 1073 624 1075
rect 311 1068 317 1070
rect 301 1065 307 1067
rect 311 1061 317 1063
rect 311 1059 313 1061
rect 315 1059 317 1061
rect 311 1057 317 1059
rect 208 1051 210 1056
rect 215 1051 217 1056
rect 222 1051 224 1056
rect 263 1051 265 1056
rect 273 1051 275 1056
rect 285 1051 287 1056
rect 295 1053 297 1056
rect 311 1053 313 1057
rect 295 1051 313 1053
rect 608 1068 610 1073
rect 621 1068 623 1073
rect 628 1068 630 1081
rect 647 1079 649 1081
rect 651 1079 658 1081
rect 666 1079 668 1086
rect 726 1110 728 1114
rect 700 1101 702 1105
rect 710 1101 712 1105
rect 737 1085 743 1087
rect 737 1083 739 1085
rect 741 1083 743 1085
rect 647 1077 658 1079
rect 656 1070 658 1077
rect 662 1077 668 1079
rect 662 1075 664 1077
rect 666 1075 668 1077
rect 662 1073 668 1075
rect 690 1080 692 1083
rect 690 1078 696 1080
rect 690 1076 692 1078
rect 694 1076 696 1078
rect 690 1074 696 1076
rect 700 1079 702 1083
rect 710 1080 712 1083
rect 726 1080 728 1083
rect 737 1081 743 1083
rect 737 1080 739 1081
rect 700 1077 706 1079
rect 710 1078 720 1080
rect 726 1078 739 1080
rect 700 1075 702 1077
rect 704 1075 706 1077
rect 663 1070 665 1073
rect 580 1056 582 1061
rect 608 1055 610 1059
rect 621 1052 623 1057
rect 628 1052 630 1057
rect 691 1065 693 1074
rect 700 1073 706 1075
rect 718 1074 720 1078
rect 700 1070 702 1073
rect 698 1068 702 1070
rect 718 1072 727 1074
rect 718 1070 723 1072
rect 725 1070 727 1072
rect 734 1070 736 1078
rect 698 1065 700 1068
rect 708 1065 710 1069
rect 718 1068 727 1070
rect 718 1065 720 1068
rect 734 1058 736 1061
rect 731 1056 736 1058
rect 656 1046 658 1050
rect 663 1046 665 1050
rect 691 1048 693 1053
rect 698 1048 700 1053
rect 708 1048 710 1056
rect 718 1052 720 1056
rect 731 1048 733 1056
rect 708 1046 733 1048
rect 90 1040 115 1042
rect 90 1032 92 1040
rect 103 1032 105 1036
rect 113 1032 115 1040
rect 123 1035 125 1040
rect 130 1035 132 1040
rect 158 1038 160 1042
rect 165 1038 167 1042
rect 87 1030 92 1032
rect 87 1027 89 1030
rect 103 1020 105 1023
rect 96 1018 105 1020
rect 113 1019 115 1023
rect 123 1020 125 1023
rect 87 1010 89 1018
rect 96 1016 98 1018
rect 100 1016 105 1018
rect 96 1014 105 1016
rect 121 1018 125 1020
rect 121 1015 123 1018
rect 103 1010 105 1014
rect 117 1013 123 1015
rect 130 1014 132 1023
rect 217 1036 219 1041
rect 227 1036 229 1041
rect 239 1036 241 1041
rect 272 1032 274 1037
rect 279 1032 281 1037
rect 286 1032 288 1037
rect 598 1038 600 1042
rect 608 1038 610 1042
rect 217 1023 219 1026
rect 227 1023 229 1026
rect 239 1023 241 1026
rect 213 1021 219 1023
rect 202 1019 208 1021
rect 158 1015 160 1018
rect 117 1011 119 1013
rect 121 1011 123 1013
rect 84 1008 97 1010
rect 103 1008 113 1010
rect 117 1009 123 1011
rect 84 1007 86 1008
rect 80 1005 86 1007
rect 95 1005 97 1008
rect 111 1005 113 1008
rect 121 1005 123 1009
rect 127 1012 133 1014
rect 127 1010 129 1012
rect 131 1010 133 1012
rect 127 1008 133 1010
rect 131 1005 133 1008
rect 155 1013 161 1015
rect 155 1011 157 1013
rect 159 1011 161 1013
rect 155 1009 161 1011
rect 165 1011 167 1018
rect 202 1017 204 1019
rect 206 1017 208 1019
rect 202 1015 208 1017
rect 192 1013 198 1015
rect 192 1011 194 1013
rect 196 1011 198 1013
rect 165 1009 176 1011
rect 192 1009 201 1011
rect 80 1003 82 1005
rect 84 1003 86 1005
rect 80 1001 86 1003
rect 111 983 113 987
rect 121 983 123 987
rect 95 974 97 978
rect 155 1002 157 1009
rect 165 1007 172 1009
rect 174 1007 176 1009
rect 165 1005 176 1007
rect 199 1006 201 1009
rect 206 1006 208 1015
rect 213 1019 215 1021
rect 217 1019 219 1021
rect 213 1017 219 1019
rect 225 1021 231 1023
rect 225 1019 227 1021
rect 229 1019 231 1021
rect 225 1017 231 1019
rect 235 1021 241 1023
rect 235 1019 237 1021
rect 239 1019 241 1021
rect 299 1028 301 1033
rect 518 1027 520 1032
rect 235 1017 241 1019
rect 213 1011 215 1017
rect 229 1012 231 1017
rect 213 1009 225 1011
rect 229 1009 232 1012
rect 213 1006 215 1009
rect 223 1006 225 1009
rect 230 1006 232 1009
rect 237 1006 239 1017
rect 272 1015 274 1019
rect 263 1013 274 1015
rect 263 1011 265 1013
rect 267 1011 269 1013
rect 263 1009 269 1011
rect 165 1002 167 1005
rect 267 1000 269 1009
rect 279 1008 281 1019
rect 286 1015 288 1019
rect 299 1015 301 1019
rect 634 1031 636 1036
rect 641 1031 643 1036
rect 722 1038 724 1042
rect 732 1038 734 1042
rect 582 1021 588 1023
rect 582 1019 584 1021
rect 586 1019 588 1021
rect 285 1013 291 1015
rect 285 1011 287 1013
rect 289 1011 291 1013
rect 285 1009 291 1011
rect 295 1013 301 1015
rect 295 1011 297 1013
rect 299 1011 301 1013
rect 295 1009 301 1011
rect 275 1006 281 1008
rect 275 1004 277 1006
rect 279 1004 281 1006
rect 275 1002 281 1004
rect 279 999 281 1002
rect 289 999 291 1009
rect 299 1004 301 1009
rect 518 1015 520 1018
rect 582 1017 588 1019
rect 518 1013 524 1015
rect 518 1011 520 1013
rect 522 1011 524 1013
rect 518 1009 524 1011
rect 518 1006 520 1009
rect 267 982 269 987
rect 586 1005 588 1017
rect 598 1015 600 1023
rect 608 1020 610 1023
rect 654 1029 656 1033
rect 680 1027 682 1032
rect 593 1013 600 1015
rect 604 1018 610 1020
rect 604 1016 606 1018
rect 608 1017 610 1018
rect 608 1016 612 1017
rect 604 1014 612 1016
rect 593 1011 595 1013
rect 597 1011 600 1013
rect 593 1010 600 1011
rect 593 1008 605 1010
rect 593 1005 595 1008
rect 603 1005 605 1008
rect 610 1005 612 1014
rect 634 1007 636 1020
rect 641 1015 643 1020
rect 654 1015 656 1020
rect 706 1021 712 1023
rect 706 1019 708 1021
rect 710 1019 712 1021
rect 640 1013 646 1015
rect 640 1011 642 1013
rect 644 1011 646 1013
rect 640 1009 646 1011
rect 650 1013 656 1015
rect 650 1011 652 1013
rect 654 1011 656 1013
rect 650 1009 656 1011
rect 630 1005 636 1007
rect 131 974 133 978
rect 155 974 157 978
rect 165 974 167 978
rect 199 974 201 978
rect 206 974 208 978
rect 213 974 215 978
rect 223 974 225 978
rect 230 974 232 978
rect 237 974 239 978
rect 279 981 281 986
rect 289 981 291 986
rect 299 981 301 986
rect 518 983 520 988
rect 630 1003 632 1005
rect 634 1003 636 1005
rect 630 1001 636 1003
rect 634 998 636 1001
rect 644 998 646 1009
rect 654 1005 656 1009
rect 680 1015 682 1018
rect 706 1017 712 1019
rect 680 1013 686 1015
rect 680 1011 682 1013
rect 684 1011 686 1013
rect 680 1009 686 1011
rect 680 1006 682 1009
rect 710 1005 712 1017
rect 722 1015 724 1023
rect 732 1020 734 1023
rect 717 1013 724 1015
rect 728 1018 734 1020
rect 728 1016 730 1018
rect 732 1017 734 1018
rect 732 1016 736 1017
rect 728 1014 736 1016
rect 717 1011 719 1013
rect 721 1011 724 1013
rect 717 1010 724 1011
rect 717 1008 729 1010
rect 717 1005 719 1008
rect 727 1005 729 1008
rect 734 1005 736 1014
rect 634 980 636 985
rect 644 980 646 985
rect 654 983 656 987
rect 680 983 682 988
rect 586 974 588 978
rect 593 974 595 978
rect 603 974 605 978
rect 610 974 612 978
rect 710 974 712 978
rect 717 974 719 978
rect 727 974 729 978
rect 734 974 736 978
rect 90 966 92 970
rect 97 966 99 970
rect 207 966 209 970
rect 123 956 125 961
rect 151 957 153 961
rect 161 959 163 964
rect 171 959 173 964
rect 90 935 92 938
rect 87 933 93 935
rect 87 931 89 933
rect 91 931 93 933
rect 87 929 93 931
rect 97 932 99 938
rect 123 935 125 938
rect 151 935 153 939
rect 161 935 163 946
rect 171 943 173 946
rect 171 941 177 943
rect 171 939 173 941
rect 175 939 177 941
rect 243 966 245 970
rect 217 957 219 961
rect 227 957 229 961
rect 518 966 520 970
rect 275 959 277 964
rect 285 959 287 964
rect 295 957 297 961
rect 275 943 277 946
rect 254 941 260 943
rect 254 939 256 941
rect 258 939 260 941
rect 171 937 177 939
rect 123 933 129 935
rect 97 930 103 932
rect 88 920 90 929
rect 97 928 99 930
rect 101 928 103 930
rect 97 926 103 928
rect 123 931 125 933
rect 127 931 129 933
rect 123 929 129 931
rect 151 933 157 935
rect 151 931 153 933
rect 155 931 157 933
rect 151 929 157 931
rect 161 933 167 935
rect 161 931 163 933
rect 165 931 167 933
rect 161 929 167 931
rect 123 926 125 929
rect 99 923 101 926
rect 151 924 153 929
rect 164 924 166 929
rect 171 924 173 937
rect 207 936 209 939
rect 207 934 213 936
rect 207 932 209 934
rect 211 932 213 934
rect 207 930 213 932
rect 217 935 219 939
rect 227 936 229 939
rect 243 936 245 939
rect 254 937 260 939
rect 271 941 277 943
rect 271 939 273 941
rect 275 939 277 941
rect 271 937 277 939
rect 254 936 256 937
rect 217 933 223 935
rect 227 934 237 936
rect 243 934 256 936
rect 217 931 219 933
rect 221 931 223 933
rect 88 907 90 912
rect 99 911 101 915
rect 123 912 125 917
rect 151 911 153 915
rect 208 921 210 930
rect 217 929 223 931
rect 235 930 237 934
rect 217 926 219 929
rect 215 924 219 926
rect 235 928 244 930
rect 235 926 240 928
rect 242 926 244 928
rect 251 926 253 934
rect 215 921 217 924
rect 225 921 227 925
rect 235 924 244 926
rect 235 921 237 924
rect 164 908 166 913
rect 171 908 173 913
rect 275 924 277 937
rect 285 935 287 946
rect 554 966 556 970
rect 528 957 530 961
rect 538 957 540 961
rect 690 966 692 970
rect 586 957 588 961
rect 596 959 598 964
rect 606 959 608 964
rect 565 941 571 943
rect 565 939 567 941
rect 569 939 571 941
rect 631 957 633 961
rect 641 957 643 962
rect 651 957 653 962
rect 661 957 663 962
rect 295 935 297 939
rect 281 933 287 935
rect 281 931 283 933
rect 285 931 287 933
rect 281 929 287 931
rect 291 933 297 935
rect 291 931 293 933
rect 295 931 297 933
rect 291 929 297 931
rect 518 936 520 939
rect 518 934 524 936
rect 518 932 520 934
rect 522 932 524 934
rect 518 930 524 932
rect 528 935 530 939
rect 538 936 540 939
rect 554 936 556 939
rect 565 937 571 939
rect 565 936 567 937
rect 528 933 534 935
rect 538 934 548 936
rect 554 934 567 936
rect 586 935 588 939
rect 596 935 598 946
rect 606 943 608 946
rect 606 941 612 943
rect 606 939 608 941
rect 610 939 612 941
rect 726 966 728 970
rect 700 957 702 961
rect 710 957 712 961
rect 737 941 743 943
rect 737 939 739 941
rect 741 939 743 941
rect 606 937 612 939
rect 528 931 530 933
rect 532 931 534 933
rect 282 924 284 929
rect 295 924 297 929
rect 251 914 253 917
rect 248 912 253 914
rect 519 921 521 930
rect 528 929 534 931
rect 546 930 548 934
rect 528 926 530 929
rect 526 924 530 926
rect 546 928 555 930
rect 546 926 551 928
rect 553 926 555 928
rect 562 926 564 934
rect 586 933 592 935
rect 586 931 588 933
rect 590 931 592 933
rect 586 929 592 931
rect 596 933 602 935
rect 596 931 598 933
rect 600 931 602 933
rect 596 929 602 931
rect 526 921 528 924
rect 536 921 538 925
rect 546 924 555 926
rect 546 921 548 924
rect 208 904 210 909
rect 215 904 217 909
rect 225 904 227 912
rect 235 908 237 912
rect 248 904 250 912
rect 225 902 250 904
rect 275 908 277 913
rect 282 908 284 913
rect 295 911 297 915
rect 586 924 588 929
rect 599 924 601 929
rect 606 924 608 937
rect 631 935 633 939
rect 641 935 643 939
rect 630 933 643 935
rect 630 931 632 933
rect 634 931 643 933
rect 630 929 643 931
rect 630 926 632 929
rect 641 926 643 929
rect 651 935 653 939
rect 661 935 663 939
rect 690 936 692 939
rect 651 933 668 935
rect 651 931 664 933
rect 666 931 668 933
rect 651 929 668 931
rect 690 934 696 936
rect 690 932 692 934
rect 694 932 696 934
rect 690 930 696 932
rect 700 935 702 939
rect 710 936 712 939
rect 726 936 728 939
rect 737 937 743 939
rect 737 936 739 937
rect 700 933 706 935
rect 710 934 720 936
rect 726 934 739 936
rect 700 931 702 933
rect 704 931 706 933
rect 651 926 653 929
rect 661 926 663 929
rect 562 914 564 917
rect 559 912 564 914
rect 519 904 521 909
rect 526 904 528 909
rect 536 904 538 912
rect 546 908 548 912
rect 559 904 561 912
rect 586 911 588 915
rect 536 902 561 904
rect 599 908 601 913
rect 606 908 608 913
rect 630 911 632 915
rect 691 921 693 930
rect 700 929 706 931
rect 718 930 720 934
rect 700 926 702 929
rect 698 924 702 926
rect 718 928 727 930
rect 718 926 723 928
rect 725 926 727 928
rect 734 926 736 934
rect 698 921 700 924
rect 708 921 710 925
rect 718 924 727 926
rect 718 921 720 924
rect 641 902 643 907
rect 651 906 653 911
rect 661 906 663 911
rect 734 914 736 917
rect 731 912 736 914
rect 691 904 693 909
rect 698 904 700 909
rect 708 904 710 912
rect 718 908 720 912
rect 731 904 733 912
rect 708 902 733 904
rect 93 893 95 898
rect 100 893 102 898
rect 123 885 125 889
rect 136 887 138 892
rect 143 887 145 892
rect 93 878 95 881
rect 85 876 95 878
rect 85 874 87 876
rect 89 874 91 876
rect 85 872 91 874
rect 89 857 91 872
rect 100 871 102 881
rect 172 885 174 889
rect 185 887 187 892
rect 192 887 194 892
rect 225 887 227 892
rect 232 887 234 892
rect 245 885 247 889
rect 271 883 273 888
rect 299 885 301 889
rect 312 887 314 892
rect 319 887 321 892
rect 96 869 102 871
rect 96 867 98 869
rect 100 867 102 869
rect 96 865 102 867
rect 123 871 125 876
rect 136 871 138 876
rect 123 869 129 871
rect 123 867 125 869
rect 127 867 129 869
rect 123 865 129 867
rect 133 869 139 871
rect 133 867 135 869
rect 137 867 139 869
rect 133 865 139 867
rect 99 857 101 865
rect 123 861 125 865
rect 133 854 135 865
rect 143 863 145 876
rect 172 871 174 876
rect 185 871 187 876
rect 172 869 178 871
rect 172 867 174 869
rect 176 867 178 869
rect 172 865 178 867
rect 182 869 188 871
rect 182 867 184 869
rect 186 867 188 869
rect 182 865 188 867
rect 143 861 149 863
rect 172 861 174 865
rect 143 859 145 861
rect 147 859 149 861
rect 143 857 149 859
rect 143 854 145 857
rect 89 839 91 843
rect 99 838 101 843
rect 123 839 125 843
rect 182 854 184 865
rect 192 863 194 876
rect 225 863 227 876
rect 232 871 234 876
rect 245 871 247 876
rect 343 884 345 889
rect 356 888 358 893
rect 363 888 365 893
rect 370 888 372 893
rect 231 869 237 871
rect 231 867 233 869
rect 235 867 237 869
rect 231 865 237 867
rect 241 869 247 871
rect 241 867 243 869
rect 245 867 247 869
rect 241 865 247 867
rect 192 861 198 863
rect 192 859 194 861
rect 196 859 198 861
rect 192 857 198 859
rect 221 861 227 863
rect 221 859 223 861
rect 225 859 227 861
rect 221 857 227 859
rect 192 854 194 857
rect 225 854 227 857
rect 235 854 237 865
rect 245 861 247 865
rect 271 871 273 874
rect 299 871 301 876
rect 312 871 314 876
rect 271 869 277 871
rect 271 867 273 869
rect 275 867 277 869
rect 271 865 277 867
rect 299 869 305 871
rect 299 867 301 869
rect 303 867 305 869
rect 299 865 305 867
rect 309 869 315 871
rect 309 867 311 869
rect 313 867 315 869
rect 309 865 315 867
rect 271 862 273 865
rect 133 836 135 841
rect 143 836 145 841
rect 172 839 174 843
rect 299 861 301 865
rect 182 836 184 841
rect 192 836 194 841
rect 225 836 227 841
rect 235 836 237 841
rect 245 839 247 843
rect 271 839 273 844
rect 309 854 311 865
rect 319 863 321 876
rect 493 887 495 892
rect 500 887 502 892
rect 513 885 515 889
rect 538 883 540 888
rect 566 887 568 892
rect 573 887 575 892
rect 343 871 345 875
rect 356 871 358 875
rect 343 869 349 871
rect 343 867 345 869
rect 347 867 349 869
rect 343 865 349 867
rect 353 869 359 871
rect 353 867 355 869
rect 357 867 359 869
rect 353 865 359 867
rect 319 861 325 863
rect 319 859 321 861
rect 323 859 325 861
rect 343 860 345 865
rect 319 857 325 859
rect 319 854 321 857
rect 299 839 301 843
rect 353 855 355 865
rect 363 864 365 875
rect 370 871 372 875
rect 370 869 381 871
rect 375 867 377 869
rect 379 867 381 869
rect 375 865 381 867
rect 363 862 369 864
rect 363 860 365 862
rect 367 860 369 862
rect 363 858 369 860
rect 363 855 365 858
rect 375 856 377 865
rect 493 863 495 876
rect 500 871 502 876
rect 513 871 515 876
rect 586 885 588 889
rect 614 885 616 889
rect 627 887 629 892
rect 634 887 636 892
rect 663 888 665 893
rect 670 888 672 893
rect 677 888 679 893
rect 717 894 719 898
rect 724 894 726 898
rect 731 894 733 898
rect 499 869 505 871
rect 499 867 501 869
rect 503 867 505 869
rect 499 865 505 867
rect 509 869 515 871
rect 509 867 511 869
rect 513 867 515 869
rect 509 865 515 867
rect 489 861 495 863
rect 489 859 491 861
rect 493 859 495 861
rect 489 857 495 859
rect 493 854 495 857
rect 503 854 505 865
rect 513 861 515 865
rect 538 871 540 874
rect 538 869 544 871
rect 538 867 540 869
rect 542 867 544 869
rect 538 865 544 867
rect 538 862 540 865
rect 566 863 568 876
rect 573 871 575 876
rect 586 871 588 876
rect 572 869 578 871
rect 572 867 574 869
rect 576 867 578 869
rect 572 865 578 867
rect 582 869 588 871
rect 582 867 584 869
rect 586 867 588 869
rect 582 865 588 867
rect 309 836 311 841
rect 319 836 321 841
rect 343 837 345 842
rect 353 837 355 842
rect 363 837 365 842
rect 375 838 377 843
rect 562 861 568 863
rect 562 859 564 861
rect 566 859 568 861
rect 562 857 568 859
rect 566 854 568 857
rect 576 854 578 865
rect 586 861 588 865
rect 614 871 616 876
rect 627 871 629 876
rect 614 869 620 871
rect 614 867 616 869
rect 618 867 620 869
rect 614 865 620 867
rect 624 869 630 871
rect 624 867 626 869
rect 628 867 630 869
rect 624 865 630 867
rect 614 861 616 865
rect 493 836 495 841
rect 503 836 505 841
rect 513 839 515 843
rect 538 839 540 844
rect 624 854 626 865
rect 634 863 636 876
rect 690 884 692 889
rect 663 871 665 875
rect 654 869 665 871
rect 654 867 656 869
rect 658 867 660 869
rect 654 865 660 867
rect 634 861 640 863
rect 634 859 636 861
rect 638 859 640 861
rect 634 857 640 859
rect 634 854 636 857
rect 658 856 660 865
rect 670 864 672 875
rect 677 871 679 875
rect 690 871 692 875
rect 717 871 719 874
rect 676 869 682 871
rect 676 867 678 869
rect 680 867 682 869
rect 676 865 682 867
rect 686 869 692 871
rect 686 867 688 869
rect 690 867 692 869
rect 686 865 692 867
rect 710 869 719 871
rect 710 867 712 869
rect 714 867 716 869
rect 710 865 716 867
rect 666 862 672 864
rect 666 860 668 862
rect 670 860 672 862
rect 666 858 672 860
rect 566 836 568 841
rect 576 836 578 841
rect 586 839 588 843
rect 614 839 616 843
rect 670 855 672 858
rect 680 855 682 865
rect 690 860 692 865
rect 624 836 626 841
rect 634 836 636 841
rect 658 838 660 843
rect 714 854 716 865
rect 724 863 726 874
rect 731 871 733 874
rect 730 869 736 871
rect 730 867 732 869
rect 734 867 736 869
rect 730 865 736 867
rect 720 861 726 863
rect 720 859 722 861
rect 724 859 726 861
rect 720 857 726 859
rect 724 854 726 857
rect 734 854 736 865
rect 670 837 672 842
rect 680 837 682 842
rect 690 837 692 842
rect 714 830 716 834
rect 724 830 726 834
rect 734 830 736 834
rect 87 822 89 826
rect 97 822 99 826
rect 107 822 109 826
rect 131 814 133 819
rect 141 814 143 819
rect 151 814 153 819
rect 87 791 89 802
rect 97 799 99 802
rect 97 797 103 799
rect 97 795 99 797
rect 101 795 103 797
rect 97 793 103 795
rect 87 789 93 791
rect 87 787 89 789
rect 91 787 93 789
rect 87 785 93 787
rect 90 782 92 785
rect 97 782 99 793
rect 107 791 109 802
rect 163 813 165 818
rect 187 815 189 820
rect 197 815 199 820
rect 131 791 133 796
rect 141 791 143 801
rect 151 798 153 801
rect 207 813 209 817
rect 235 813 237 817
rect 245 815 247 820
rect 255 815 257 820
rect 151 796 157 798
rect 151 794 153 796
rect 155 794 157 796
rect 151 792 157 794
rect 107 789 113 791
rect 107 787 109 789
rect 111 787 113 789
rect 104 785 113 787
rect 131 789 137 791
rect 131 787 133 789
rect 135 787 137 789
rect 131 785 137 787
rect 141 789 147 791
rect 141 787 143 789
rect 145 787 147 789
rect 141 785 147 787
rect 104 782 106 785
rect 131 781 133 785
rect 144 781 146 785
rect 151 781 153 792
rect 163 791 165 800
rect 187 799 189 802
rect 183 797 189 799
rect 183 795 185 797
rect 187 795 189 797
rect 183 793 189 795
rect 163 789 169 791
rect 163 787 165 789
rect 167 787 169 789
rect 158 785 169 787
rect 158 781 160 785
rect 131 767 133 772
rect 187 780 189 793
rect 197 791 199 802
rect 283 812 285 817
rect 308 813 310 817
rect 318 815 320 820
rect 328 815 330 820
rect 207 791 209 795
rect 193 789 199 791
rect 193 787 195 789
rect 197 787 199 789
rect 193 785 199 787
rect 203 789 209 791
rect 203 787 205 789
rect 207 787 209 789
rect 203 785 209 787
rect 194 780 196 785
rect 207 780 209 785
rect 235 791 237 795
rect 245 791 247 802
rect 255 799 257 802
rect 255 797 261 799
rect 255 795 257 797
rect 259 795 261 797
rect 255 793 261 795
rect 446 813 448 818
rect 458 814 460 819
rect 468 814 470 819
rect 478 814 480 819
rect 502 815 504 820
rect 512 815 514 820
rect 235 789 241 791
rect 235 787 237 789
rect 239 787 241 789
rect 235 785 241 787
rect 245 789 251 791
rect 245 787 247 789
rect 249 787 251 789
rect 245 785 251 787
rect 235 780 237 785
rect 248 780 250 785
rect 255 780 257 793
rect 283 791 285 794
rect 279 789 285 791
rect 279 787 281 789
rect 283 787 285 789
rect 279 785 285 787
rect 283 782 285 785
rect 308 791 310 795
rect 318 791 320 802
rect 328 799 330 802
rect 328 797 334 799
rect 328 795 330 797
rect 332 795 334 797
rect 328 793 334 795
rect 308 789 314 791
rect 308 787 310 789
rect 312 787 314 789
rect 308 785 314 787
rect 318 789 324 791
rect 318 787 320 789
rect 322 787 324 789
rect 318 785 324 787
rect 90 758 92 762
rect 97 758 99 762
rect 104 758 106 762
rect 144 763 146 768
rect 151 763 153 768
rect 158 763 160 768
rect 187 764 189 769
rect 194 764 196 769
rect 207 767 209 771
rect 235 767 237 771
rect 308 780 310 785
rect 321 780 323 785
rect 328 780 330 793
rect 446 791 448 800
rect 458 798 460 801
rect 454 796 460 798
rect 454 794 456 796
rect 458 794 460 796
rect 454 792 460 794
rect 442 789 448 791
rect 442 787 444 789
rect 446 787 448 789
rect 442 785 453 787
rect 451 781 453 785
rect 458 781 460 792
rect 468 791 470 801
rect 522 813 524 817
rect 502 799 504 802
rect 498 797 504 799
rect 478 791 480 796
rect 498 795 500 797
rect 502 795 504 797
rect 498 793 504 795
rect 464 789 470 791
rect 464 787 466 789
rect 468 787 470 789
rect 464 785 470 787
rect 474 789 480 791
rect 474 787 476 789
rect 478 787 480 789
rect 474 785 480 787
rect 465 781 467 785
rect 478 781 480 785
rect 248 764 250 769
rect 255 764 257 769
rect 283 768 285 773
rect 308 767 310 771
rect 321 764 323 769
rect 328 764 330 769
rect 502 780 504 793
rect 512 791 514 802
rect 550 812 552 817
rect 576 813 578 817
rect 586 815 588 820
rect 596 815 598 820
rect 629 815 631 820
rect 639 815 641 820
rect 522 791 524 795
rect 649 813 651 817
rect 678 815 680 820
rect 688 815 690 820
rect 550 791 552 794
rect 508 789 514 791
rect 508 787 510 789
rect 512 787 514 789
rect 508 785 514 787
rect 518 789 524 791
rect 518 787 520 789
rect 522 787 524 789
rect 518 785 524 787
rect 546 789 552 791
rect 546 787 548 789
rect 550 787 552 789
rect 546 785 552 787
rect 509 780 511 785
rect 522 780 524 785
rect 550 782 552 785
rect 576 791 578 795
rect 586 791 588 802
rect 596 799 598 802
rect 629 799 631 802
rect 596 797 602 799
rect 596 795 598 797
rect 600 795 602 797
rect 596 793 602 795
rect 625 797 631 799
rect 625 795 627 797
rect 629 795 631 797
rect 625 793 631 795
rect 576 789 582 791
rect 576 787 578 789
rect 580 787 582 789
rect 576 785 582 787
rect 586 789 592 791
rect 586 787 588 789
rect 590 787 592 789
rect 586 785 592 787
rect 451 763 453 768
rect 458 763 460 768
rect 465 763 467 768
rect 478 767 480 772
rect 576 780 578 785
rect 589 780 591 785
rect 596 780 598 793
rect 629 780 631 793
rect 639 791 641 802
rect 698 813 700 817
rect 722 813 724 818
rect 732 813 734 817
rect 678 799 680 802
rect 674 797 680 799
rect 674 795 676 797
rect 678 795 680 797
rect 649 791 651 795
rect 674 793 680 795
rect 635 789 641 791
rect 635 787 637 789
rect 639 787 641 789
rect 635 785 641 787
rect 645 789 651 791
rect 645 787 647 789
rect 649 787 651 789
rect 645 785 651 787
rect 636 780 638 785
rect 649 780 651 785
rect 678 780 680 793
rect 688 791 690 802
rect 698 791 700 795
rect 722 791 724 799
rect 684 789 690 791
rect 684 787 686 789
rect 688 787 690 789
rect 684 785 690 787
rect 694 789 700 791
rect 694 787 696 789
rect 698 787 700 789
rect 694 785 700 787
rect 685 780 687 785
rect 698 780 700 785
rect 721 789 727 791
rect 721 787 723 789
rect 725 787 727 789
rect 721 785 727 787
rect 502 764 504 769
rect 509 764 511 769
rect 522 767 524 771
rect 550 768 552 773
rect 576 767 578 771
rect 589 764 591 769
rect 596 764 598 769
rect 629 764 631 769
rect 636 764 638 769
rect 649 767 651 771
rect 721 775 723 785
rect 732 784 734 799
rect 732 782 738 784
rect 732 780 734 782
rect 736 780 738 782
rect 728 778 738 780
rect 728 775 730 778
rect 678 764 680 769
rect 685 764 687 769
rect 698 767 700 771
rect 721 758 723 763
rect 728 758 730 763
rect 90 752 115 754
rect 90 744 92 752
rect 103 744 105 748
rect 113 744 115 752
rect 123 747 125 752
rect 130 747 132 752
rect 87 742 92 744
rect 87 739 89 742
rect 160 745 162 750
rect 170 745 172 750
rect 180 749 182 754
rect 103 732 105 735
rect 96 730 105 732
rect 113 731 115 735
rect 123 732 125 735
rect 87 722 89 730
rect 96 728 98 730
rect 100 728 105 730
rect 96 726 105 728
rect 121 730 125 732
rect 121 727 123 730
rect 103 722 105 726
rect 117 725 123 727
rect 130 726 132 735
rect 191 741 193 745
rect 215 743 217 748
rect 222 743 224 748
rect 262 752 287 754
rect 235 741 237 745
rect 262 744 264 752
rect 275 744 277 748
rect 285 744 287 752
rect 295 747 297 752
rect 302 747 304 752
rect 259 742 264 744
rect 259 739 261 742
rect 160 727 162 730
rect 170 727 172 730
rect 117 723 119 725
rect 121 723 123 725
rect 84 720 97 722
rect 103 720 113 722
rect 117 721 123 723
rect 84 719 86 720
rect 80 717 86 719
rect 95 717 97 720
rect 111 717 113 720
rect 121 717 123 721
rect 127 724 133 726
rect 127 722 129 724
rect 131 722 133 724
rect 127 720 133 722
rect 155 725 172 727
rect 155 723 157 725
rect 159 723 172 725
rect 155 721 172 723
rect 131 717 133 720
rect 160 717 162 721
rect 170 717 172 721
rect 180 727 182 730
rect 191 727 193 730
rect 180 725 193 727
rect 180 723 189 725
rect 191 723 193 725
rect 180 721 193 723
rect 180 717 182 721
rect 190 717 192 721
rect 215 719 217 732
rect 222 727 224 732
rect 235 727 237 732
rect 327 739 329 744
rect 526 741 528 745
rect 539 743 541 748
rect 546 743 548 748
rect 573 752 598 754
rect 573 744 575 752
rect 586 744 588 748
rect 596 744 598 752
rect 606 747 608 752
rect 613 747 615 752
rect 275 732 277 735
rect 268 730 277 732
rect 285 731 287 735
rect 295 732 297 735
rect 221 725 227 727
rect 221 723 223 725
rect 225 723 227 725
rect 221 721 227 723
rect 231 725 237 727
rect 231 723 233 725
rect 235 723 237 725
rect 231 721 237 723
rect 259 722 261 730
rect 268 728 270 730
rect 272 728 277 730
rect 268 726 277 728
rect 293 730 297 732
rect 293 727 295 730
rect 275 722 277 726
rect 289 725 295 727
rect 302 726 304 735
rect 570 742 575 744
rect 570 739 572 742
rect 327 727 329 730
rect 526 727 528 732
rect 539 727 541 732
rect 289 723 291 725
rect 293 723 295 725
rect 211 717 217 719
rect 80 715 82 717
rect 84 715 86 717
rect 80 713 86 715
rect 111 695 113 699
rect 121 695 123 699
rect 95 686 97 690
rect 211 715 213 717
rect 215 715 217 717
rect 211 713 217 715
rect 215 710 217 713
rect 225 710 227 721
rect 235 717 237 721
rect 256 720 269 722
rect 275 720 285 722
rect 289 721 295 723
rect 256 719 258 720
rect 252 717 258 719
rect 267 717 269 720
rect 283 717 285 720
rect 293 717 295 721
rect 299 724 305 726
rect 299 722 301 724
rect 303 722 305 724
rect 299 720 305 722
rect 303 717 305 720
rect 327 725 333 727
rect 327 723 329 725
rect 331 723 333 725
rect 327 721 333 723
rect 526 725 532 727
rect 526 723 528 725
rect 530 723 532 725
rect 526 721 532 723
rect 536 725 542 727
rect 536 723 538 725
rect 540 723 542 725
rect 536 721 542 723
rect 327 718 329 721
rect 160 694 162 699
rect 170 694 172 699
rect 180 694 182 699
rect 190 695 192 699
rect 252 715 254 717
rect 256 715 258 717
rect 252 713 258 715
rect 215 692 217 697
rect 225 692 227 697
rect 235 695 237 699
rect 131 686 133 690
rect 283 695 285 699
rect 293 695 295 699
rect 267 686 269 690
rect 526 717 528 721
rect 327 695 329 700
rect 536 710 538 721
rect 546 719 548 732
rect 650 743 652 748
rect 657 743 659 748
rect 586 732 588 735
rect 579 730 588 732
rect 596 731 598 735
rect 606 732 608 735
rect 570 722 572 730
rect 579 728 581 730
rect 583 728 588 730
rect 579 726 588 728
rect 604 730 608 732
rect 604 727 606 730
rect 586 722 588 726
rect 600 725 606 727
rect 613 726 615 735
rect 670 741 672 745
rect 698 739 700 744
rect 722 741 724 745
rect 733 744 735 749
rect 600 723 602 725
rect 604 723 606 725
rect 567 720 580 722
rect 586 720 596 722
rect 600 721 606 723
rect 567 719 569 720
rect 546 717 552 719
rect 546 715 548 717
rect 550 715 552 717
rect 546 713 552 715
rect 563 717 569 719
rect 578 717 580 720
rect 594 717 596 720
rect 604 717 606 721
rect 610 724 616 726
rect 610 722 612 724
rect 614 722 616 724
rect 610 720 616 722
rect 614 717 616 720
rect 650 719 652 732
rect 657 727 659 732
rect 670 727 672 732
rect 722 730 724 733
rect 698 727 700 730
rect 656 725 662 727
rect 656 723 658 725
rect 660 723 662 725
rect 656 721 662 723
rect 666 725 672 727
rect 666 723 668 725
rect 670 723 672 725
rect 666 721 672 723
rect 694 725 700 727
rect 694 723 696 725
rect 698 723 700 725
rect 720 728 726 730
rect 720 726 722 728
rect 724 726 726 728
rect 733 727 735 736
rect 720 724 726 726
rect 694 721 700 723
rect 646 717 652 719
rect 563 715 565 717
rect 567 715 569 717
rect 563 713 569 715
rect 546 710 548 713
rect 526 695 528 699
rect 303 686 305 690
rect 536 692 538 697
rect 546 692 548 697
rect 594 695 596 699
rect 604 695 606 699
rect 578 686 580 690
rect 646 715 648 717
rect 650 715 652 717
rect 646 713 652 715
rect 650 710 652 713
rect 660 710 662 721
rect 670 717 672 721
rect 698 718 700 721
rect 724 718 726 724
rect 730 725 736 727
rect 730 723 732 725
rect 734 723 736 725
rect 730 721 736 723
rect 731 718 733 721
rect 650 692 652 697
rect 660 692 662 697
rect 670 695 672 699
rect 698 695 700 700
rect 614 686 616 690
rect 724 686 726 690
rect 731 686 733 690
rect 87 678 89 682
rect 94 678 96 682
rect 104 678 106 682
rect 111 678 113 682
rect 211 678 213 682
rect 218 678 220 682
rect 228 678 230 682
rect 235 678 237 682
rect 141 668 143 673
rect 167 669 169 673
rect 177 671 179 676
rect 187 671 189 676
rect 87 642 89 651
rect 94 648 96 651
rect 104 648 106 651
rect 94 646 106 648
rect 99 645 106 646
rect 99 643 102 645
rect 104 643 106 645
rect 87 640 95 642
rect 87 639 91 640
rect 89 638 91 639
rect 93 638 95 640
rect 89 636 95 638
rect 99 641 106 643
rect 89 633 91 636
rect 99 633 101 641
rect 111 639 113 651
rect 141 647 143 650
rect 137 645 143 647
rect 137 643 139 645
rect 141 643 143 645
rect 137 641 143 643
rect 111 637 117 639
rect 141 638 143 641
rect 167 647 169 651
rect 177 647 179 658
rect 187 655 189 658
rect 187 653 193 655
rect 187 651 189 653
rect 191 651 193 653
rect 522 670 524 675
rect 532 670 534 675
rect 542 670 544 675
rect 584 678 586 682
rect 591 678 593 682
rect 598 678 600 682
rect 608 678 610 682
rect 615 678 617 682
rect 622 678 624 682
rect 656 678 658 682
rect 666 678 668 682
rect 690 678 692 682
rect 554 669 556 674
rect 187 649 193 651
rect 167 645 173 647
rect 167 643 169 645
rect 171 643 173 645
rect 167 641 173 643
rect 177 645 183 647
rect 177 643 179 645
rect 181 643 183 645
rect 177 641 183 643
rect 111 635 113 637
rect 115 635 117 637
rect 111 633 117 635
rect 167 636 169 641
rect 180 636 182 641
rect 187 636 189 649
rect 211 642 213 651
rect 218 648 220 651
rect 228 648 230 651
rect 218 646 230 648
rect 223 645 230 646
rect 223 643 226 645
rect 228 643 230 645
rect 211 640 219 642
rect 211 639 215 640
rect 213 638 215 639
rect 217 638 219 640
rect 213 636 219 638
rect 223 641 230 643
rect 141 624 143 629
rect 167 623 169 627
rect 213 633 215 636
rect 223 633 225 641
rect 235 639 237 651
rect 522 647 524 652
rect 532 647 534 657
rect 542 654 544 657
rect 542 652 548 654
rect 542 650 544 652
rect 546 650 548 652
rect 542 648 548 650
rect 522 645 528 647
rect 522 643 524 645
rect 526 643 528 645
rect 522 641 528 643
rect 532 645 538 647
rect 532 643 534 645
rect 536 643 538 645
rect 532 641 538 643
rect 235 637 241 639
rect 522 637 524 641
rect 535 637 537 641
rect 542 637 544 648
rect 554 647 556 656
rect 656 651 658 654
rect 554 645 560 647
rect 554 643 556 645
rect 558 643 560 645
rect 549 641 560 643
rect 549 637 551 641
rect 584 639 586 650
rect 591 647 593 650
rect 598 647 600 650
rect 608 647 610 650
rect 591 644 594 647
rect 598 645 610 647
rect 592 639 594 644
rect 608 639 610 645
rect 582 637 588 639
rect 235 635 237 637
rect 239 635 241 637
rect 235 633 241 635
rect 89 614 91 618
rect 99 614 101 618
rect 180 620 182 625
rect 187 620 189 625
rect 522 623 524 628
rect 582 635 584 637
rect 586 635 588 637
rect 582 633 588 635
rect 592 637 598 639
rect 592 635 594 637
rect 596 635 598 637
rect 592 633 598 635
rect 604 637 610 639
rect 604 635 606 637
rect 608 635 610 637
rect 615 641 617 650
rect 622 647 624 650
rect 647 649 658 651
rect 647 647 649 649
rect 651 647 658 649
rect 666 647 668 654
rect 726 678 728 682
rect 700 669 702 673
rect 710 669 712 673
rect 737 653 743 655
rect 737 651 739 653
rect 741 651 743 653
rect 622 645 631 647
rect 647 645 658 647
rect 625 643 627 645
rect 629 643 631 645
rect 625 641 631 643
rect 615 639 621 641
rect 615 637 617 639
rect 619 637 621 639
rect 656 638 658 645
rect 662 645 668 647
rect 662 643 664 645
rect 666 643 668 645
rect 662 641 668 643
rect 690 648 692 651
rect 690 646 696 648
rect 690 644 692 646
rect 694 644 696 646
rect 690 642 696 644
rect 700 647 702 651
rect 710 648 712 651
rect 726 648 728 651
rect 737 649 743 651
rect 737 648 739 649
rect 700 645 706 647
rect 710 646 720 648
rect 726 646 739 648
rect 700 643 702 645
rect 704 643 706 645
rect 663 638 665 641
rect 615 635 621 637
rect 604 633 610 635
rect 582 630 584 633
rect 594 630 596 633
rect 604 630 606 633
rect 213 614 215 618
rect 223 614 225 618
rect 535 619 537 624
rect 542 619 544 624
rect 549 619 551 624
rect 582 615 584 620
rect 594 615 596 620
rect 604 615 606 620
rect 691 633 693 642
rect 700 641 706 643
rect 718 642 720 646
rect 700 638 702 641
rect 698 636 702 638
rect 718 640 727 642
rect 718 638 723 640
rect 725 638 727 640
rect 734 638 736 646
rect 698 633 700 636
rect 708 633 710 637
rect 718 636 727 638
rect 718 633 720 636
rect 734 626 736 629
rect 731 624 736 626
rect 656 614 658 618
rect 663 614 665 618
rect 691 616 693 621
rect 698 616 700 621
rect 708 616 710 624
rect 718 620 720 624
rect 731 616 733 624
rect 708 614 733 616
rect 90 608 115 610
rect 90 600 92 608
rect 103 600 105 604
rect 113 600 115 608
rect 123 603 125 608
rect 130 603 132 608
rect 158 606 160 610
rect 165 606 167 610
rect 87 598 92 600
rect 87 595 89 598
rect 103 588 105 591
rect 96 586 105 588
rect 113 587 115 591
rect 123 588 125 591
rect 87 578 89 586
rect 96 584 98 586
rect 100 584 105 586
rect 96 582 105 584
rect 121 586 125 588
rect 121 583 123 586
rect 103 578 105 582
rect 117 581 123 583
rect 130 582 132 591
rect 193 599 195 604
rect 200 599 202 604
rect 213 597 215 601
rect 241 595 243 600
rect 158 583 160 586
rect 117 579 119 581
rect 121 579 123 581
rect 84 576 97 578
rect 103 576 113 578
rect 117 577 123 579
rect 84 575 86 576
rect 80 573 86 575
rect 95 573 97 576
rect 111 573 113 576
rect 121 573 123 577
rect 127 580 133 582
rect 127 578 129 580
rect 131 578 133 580
rect 127 576 133 578
rect 131 573 133 576
rect 155 581 161 583
rect 155 579 157 581
rect 159 579 161 581
rect 155 577 161 579
rect 165 579 167 586
rect 165 577 176 579
rect 80 571 82 573
rect 84 571 86 573
rect 80 569 86 571
rect 111 551 113 555
rect 121 551 123 555
rect 95 542 97 546
rect 155 570 157 577
rect 165 575 172 577
rect 174 575 176 577
rect 193 575 195 588
rect 200 583 202 588
rect 213 583 215 588
rect 510 603 528 605
rect 510 599 512 603
rect 526 600 528 603
rect 536 600 538 605
rect 548 600 550 605
rect 558 600 560 605
rect 599 600 601 605
rect 606 600 608 605
rect 613 600 615 605
rect 506 597 512 599
rect 506 595 508 597
rect 510 595 512 597
rect 506 593 512 595
rect 516 589 522 591
rect 506 586 512 588
rect 199 581 205 583
rect 199 579 201 581
rect 203 579 205 581
rect 199 577 205 579
rect 209 581 215 583
rect 209 579 211 581
rect 213 579 215 581
rect 209 577 215 579
rect 165 573 176 575
rect 189 573 195 575
rect 165 570 167 573
rect 189 571 191 573
rect 193 571 195 573
rect 189 569 195 571
rect 193 566 195 569
rect 203 566 205 577
rect 213 573 215 577
rect 241 583 243 586
rect 506 584 508 586
rect 510 584 512 586
rect 241 581 247 583
rect 506 582 512 584
rect 516 587 518 589
rect 520 587 522 589
rect 516 585 522 587
rect 241 579 243 581
rect 245 579 247 581
rect 241 577 247 579
rect 496 580 502 582
rect 496 578 498 580
rect 500 578 502 580
rect 241 574 243 577
rect 496 576 504 578
rect 502 573 504 576
rect 509 573 511 582
rect 516 573 518 585
rect 526 578 528 594
rect 536 591 538 594
rect 535 589 541 591
rect 548 589 550 594
rect 535 587 537 589
rect 539 587 541 589
rect 535 585 541 587
rect 539 579 541 585
rect 546 587 552 589
rect 546 585 548 587
rect 550 585 552 587
rect 546 583 552 585
rect 523 576 535 578
rect 539 576 542 579
rect 523 573 525 576
rect 533 573 535 576
rect 540 573 542 576
rect 547 573 549 583
rect 558 582 560 594
rect 626 596 628 601
rect 650 599 652 604
rect 657 599 659 604
rect 724 606 726 610
rect 731 606 733 610
rect 670 597 672 601
rect 698 595 700 600
rect 599 583 601 587
rect 558 580 567 582
rect 558 578 563 580
rect 565 578 567 580
rect 554 576 567 578
rect 590 581 601 583
rect 590 579 592 581
rect 594 579 596 581
rect 590 577 596 579
rect 554 573 556 576
rect 193 548 195 553
rect 203 548 205 553
rect 213 551 215 555
rect 241 551 243 556
rect 502 551 504 555
rect 509 551 511 555
rect 516 551 518 555
rect 523 551 525 555
rect 131 542 133 546
rect 155 542 157 546
rect 165 542 167 546
rect 594 568 596 577
rect 606 576 608 587
rect 613 583 615 587
rect 626 583 628 587
rect 612 581 618 583
rect 612 579 614 581
rect 616 579 618 581
rect 612 577 618 579
rect 622 581 628 583
rect 622 579 624 581
rect 626 579 628 581
rect 622 577 628 579
rect 602 574 608 576
rect 602 572 604 574
rect 606 572 608 574
rect 602 570 608 572
rect 606 567 608 570
rect 616 567 618 577
rect 626 572 628 577
rect 650 575 652 588
rect 657 583 659 588
rect 670 583 672 588
rect 698 583 700 586
rect 656 581 662 583
rect 656 579 658 581
rect 660 579 662 581
rect 656 577 662 579
rect 666 581 672 583
rect 666 579 668 581
rect 670 579 672 581
rect 666 577 672 579
rect 694 581 700 583
rect 694 579 696 581
rect 698 579 700 581
rect 724 579 726 586
rect 731 583 733 586
rect 694 577 700 579
rect 646 573 652 575
rect 594 550 596 555
rect 646 571 648 573
rect 650 571 652 573
rect 646 569 652 571
rect 650 566 652 569
rect 660 566 662 577
rect 670 573 672 577
rect 698 574 700 577
rect 715 577 726 579
rect 730 581 736 583
rect 730 579 732 581
rect 734 579 736 581
rect 730 577 736 579
rect 715 575 717 577
rect 719 575 726 577
rect 533 543 535 548
rect 540 543 542 548
rect 547 543 549 548
rect 554 543 556 548
rect 606 549 608 554
rect 616 549 618 554
rect 626 549 628 554
rect 715 573 726 575
rect 724 570 726 573
rect 734 570 736 577
rect 650 548 652 553
rect 660 548 662 553
rect 670 551 672 555
rect 698 551 700 556
rect 724 542 726 546
rect 734 542 736 546
rect 87 534 89 538
rect 94 534 96 538
rect 104 534 106 538
rect 111 534 113 538
rect 166 534 168 538
rect 139 524 141 529
rect 87 498 89 507
rect 94 504 96 507
rect 104 504 106 507
rect 94 502 106 504
rect 99 501 106 502
rect 99 499 102 501
rect 104 499 106 501
rect 87 496 95 498
rect 87 495 91 496
rect 89 494 91 495
rect 93 494 95 496
rect 89 492 95 494
rect 99 497 106 499
rect 89 489 91 492
rect 99 489 101 497
rect 111 495 113 507
rect 202 534 204 538
rect 176 525 178 529
rect 186 525 188 529
rect 247 533 249 537
rect 237 525 239 529
rect 213 509 219 511
rect 486 530 488 535
rect 496 530 498 535
rect 506 530 508 535
rect 516 530 518 535
rect 542 534 544 538
rect 456 524 458 529
rect 213 507 215 509
rect 217 507 219 509
rect 139 503 141 506
rect 135 501 141 503
rect 135 499 137 501
rect 139 499 141 501
rect 135 497 141 499
rect 166 504 168 507
rect 166 502 172 504
rect 166 500 168 502
rect 170 500 172 502
rect 166 498 172 500
rect 176 503 178 507
rect 186 504 188 507
rect 202 504 204 507
rect 213 505 219 507
rect 213 504 215 505
rect 237 504 239 509
rect 247 504 249 509
rect 176 501 182 503
rect 186 502 196 504
rect 202 502 215 504
rect 229 502 249 504
rect 456 503 458 506
rect 486 503 488 513
rect 496 510 498 513
rect 506 510 508 513
rect 492 508 498 510
rect 492 506 494 508
rect 496 506 498 508
rect 492 504 498 506
rect 502 508 508 510
rect 502 506 504 508
rect 506 506 508 508
rect 502 504 508 506
rect 176 499 178 501
rect 180 499 182 501
rect 111 493 117 495
rect 139 494 141 497
rect 111 491 113 493
rect 115 491 117 493
rect 111 489 117 491
rect 167 489 169 498
rect 176 497 182 499
rect 194 498 196 502
rect 176 494 178 497
rect 174 492 178 494
rect 194 496 203 498
rect 194 494 199 496
rect 201 494 203 496
rect 210 494 212 502
rect 229 500 231 502
rect 233 500 239 502
rect 229 498 239 500
rect 237 494 239 498
rect 247 494 249 502
rect 452 501 458 503
rect 452 499 454 501
rect 456 499 458 501
rect 452 497 458 499
rect 480 501 488 503
rect 480 499 482 501
rect 484 499 488 501
rect 480 497 491 499
rect 456 494 458 497
rect 489 494 491 497
rect 496 494 498 504
rect 503 494 505 504
rect 516 503 518 513
rect 578 534 580 538
rect 552 525 554 529
rect 562 525 564 529
rect 656 534 658 538
rect 663 534 665 538
rect 690 534 692 538
rect 610 527 612 532
rect 620 527 622 532
rect 630 525 632 529
rect 610 511 612 514
rect 589 509 595 511
rect 589 507 591 509
rect 593 507 595 509
rect 512 501 518 503
rect 512 500 514 501
rect 510 499 514 500
rect 516 499 518 501
rect 510 497 518 499
rect 542 504 544 507
rect 542 502 548 504
rect 542 500 544 502
rect 546 500 548 502
rect 542 498 548 500
rect 552 503 554 507
rect 562 504 564 507
rect 578 504 580 507
rect 589 505 595 507
rect 606 509 612 511
rect 606 507 608 509
rect 610 507 612 509
rect 606 505 612 507
rect 589 504 591 505
rect 552 501 558 503
rect 562 502 572 504
rect 578 502 591 504
rect 552 499 554 501
rect 556 499 558 501
rect 510 494 512 497
rect 174 489 176 492
rect 184 489 186 493
rect 194 492 203 494
rect 194 489 196 492
rect 139 480 141 485
rect 210 482 212 485
rect 207 480 212 482
rect 89 470 91 474
rect 99 470 101 474
rect 167 472 169 477
rect 174 472 176 477
rect 184 472 186 480
rect 194 476 196 480
rect 207 472 209 480
rect 237 479 239 484
rect 247 479 249 484
rect 456 480 458 485
rect 184 470 209 472
rect 543 489 545 498
rect 552 497 558 499
rect 570 498 572 502
rect 552 494 554 497
rect 550 492 554 494
rect 570 496 579 498
rect 570 494 575 496
rect 577 494 579 496
rect 586 494 588 502
rect 550 489 552 492
rect 560 489 562 493
rect 570 492 579 494
rect 570 489 572 492
rect 610 492 612 505
rect 620 503 622 514
rect 630 503 632 507
rect 726 534 728 538
rect 700 525 702 529
rect 710 525 712 529
rect 737 509 743 511
rect 737 507 739 509
rect 741 507 743 509
rect 616 501 622 503
rect 616 499 618 501
rect 620 499 622 501
rect 616 497 622 499
rect 626 501 632 503
rect 626 499 628 501
rect 630 499 632 501
rect 656 500 658 506
rect 663 503 665 506
rect 690 504 692 507
rect 626 497 632 499
rect 617 492 619 497
rect 630 492 632 497
rect 652 498 658 500
rect 652 496 654 498
rect 656 496 658 498
rect 662 501 668 503
rect 662 499 664 501
rect 666 499 668 501
rect 662 497 668 499
rect 690 502 696 504
rect 690 500 692 502
rect 694 500 696 502
rect 690 498 696 500
rect 700 503 702 507
rect 710 504 712 507
rect 726 504 728 507
rect 737 505 743 507
rect 737 504 739 505
rect 700 501 706 503
rect 710 502 720 504
rect 726 502 739 504
rect 700 499 702 501
rect 704 499 706 501
rect 652 494 658 496
rect 586 482 588 485
rect 583 480 588 482
rect 654 491 656 494
rect 665 488 667 497
rect 691 489 693 498
rect 700 497 706 499
rect 718 498 720 502
rect 700 494 702 497
rect 698 492 702 494
rect 718 496 727 498
rect 718 494 723 496
rect 725 494 727 496
rect 734 494 736 502
rect 698 489 700 492
rect 708 489 710 493
rect 718 492 727 494
rect 718 489 720 492
rect 489 470 491 474
rect 496 470 498 474
rect 503 470 505 474
rect 510 470 512 474
rect 543 472 545 477
rect 550 472 552 477
rect 560 472 562 480
rect 570 476 572 480
rect 583 472 585 480
rect 560 470 585 472
rect 610 476 612 481
rect 617 476 619 481
rect 630 479 632 483
rect 654 479 656 483
rect 665 475 667 480
rect 734 482 736 485
rect 731 480 736 482
rect 691 472 693 477
rect 698 472 700 477
rect 708 472 710 480
rect 718 476 720 480
rect 731 472 733 480
rect 708 470 733 472
rect 45 361 90 363
rect 45 356 47 361
rect 14 350 16 354
rect 25 351 27 356
rect 35 351 37 356
rect 55 353 57 357
rect 45 341 47 345
rect 75 352 77 357
rect 88 349 90 361
rect 145 361 190 363
rect 145 356 147 361
rect 114 350 116 354
rect 125 351 127 356
rect 135 351 137 356
rect 14 336 16 340
rect 25 336 27 340
rect 10 334 16 336
rect 10 332 12 334
rect 14 332 16 334
rect 10 330 16 332
rect 21 334 27 336
rect 35 337 37 340
rect 35 335 49 337
rect 21 332 23 334
rect 25 332 27 334
rect 21 330 27 332
rect 43 334 49 335
rect 43 332 45 334
rect 47 332 49 334
rect 12 327 14 330
rect 23 327 25 330
rect 33 327 35 331
rect 43 330 49 332
rect 55 336 57 342
rect 75 337 77 342
rect 88 339 90 342
rect 155 353 157 357
rect 145 341 147 345
rect 175 352 177 357
rect 188 349 190 361
rect 245 361 290 363
rect 245 356 247 361
rect 214 350 216 354
rect 225 351 227 356
rect 235 351 237 356
rect 84 337 90 339
rect 55 334 64 336
rect 55 332 60 334
rect 62 332 64 334
rect 55 330 64 332
rect 74 335 80 337
rect 74 333 76 335
rect 78 333 80 335
rect 84 335 86 337
rect 88 335 90 337
rect 114 336 116 340
rect 125 336 127 340
rect 84 333 90 335
rect 74 331 80 333
rect 43 327 45 330
rect 57 327 59 330
rect 75 327 77 331
rect 12 309 14 314
rect 88 319 90 333
rect 110 334 116 336
rect 110 332 112 334
rect 114 332 116 334
rect 110 330 116 332
rect 121 334 127 336
rect 135 337 137 340
rect 135 335 149 337
rect 121 332 123 334
rect 125 332 127 334
rect 121 330 127 332
rect 143 334 149 335
rect 143 332 145 334
rect 147 332 149 334
rect 112 327 114 330
rect 123 327 125 330
rect 133 327 135 331
rect 143 330 149 332
rect 155 336 157 342
rect 175 337 177 342
rect 188 339 190 342
rect 255 353 257 357
rect 245 341 247 345
rect 275 352 277 357
rect 288 349 290 361
rect 345 361 390 363
rect 345 356 347 361
rect 314 350 316 354
rect 325 351 327 356
rect 335 351 337 356
rect 184 337 190 339
rect 155 334 164 336
rect 155 332 160 334
rect 162 332 164 334
rect 155 330 164 332
rect 174 335 180 337
rect 174 333 176 335
rect 178 333 180 335
rect 184 335 186 337
rect 188 335 190 337
rect 214 336 216 340
rect 225 336 227 340
rect 184 333 190 335
rect 174 331 180 333
rect 143 327 145 330
rect 157 327 159 330
rect 175 327 177 331
rect 75 309 77 314
rect 112 309 114 314
rect 23 300 25 305
rect 33 297 35 305
rect 43 301 45 305
rect 57 301 59 305
rect 88 297 90 309
rect 188 319 190 333
rect 210 334 216 336
rect 210 332 212 334
rect 214 332 216 334
rect 210 330 216 332
rect 221 334 227 336
rect 235 337 237 340
rect 235 335 249 337
rect 221 332 223 334
rect 225 332 227 334
rect 221 330 227 332
rect 243 334 249 335
rect 243 332 245 334
rect 247 332 249 334
rect 212 327 214 330
rect 223 327 225 330
rect 233 327 235 331
rect 243 330 249 332
rect 255 336 257 342
rect 275 337 277 342
rect 288 339 290 342
rect 355 353 357 357
rect 345 341 347 345
rect 375 352 377 357
rect 388 349 390 361
rect 445 361 490 363
rect 445 356 447 361
rect 414 350 416 354
rect 425 351 427 356
rect 435 351 437 356
rect 284 337 290 339
rect 255 334 264 336
rect 255 332 260 334
rect 262 332 264 334
rect 255 330 264 332
rect 274 335 280 337
rect 274 333 276 335
rect 278 333 280 335
rect 284 335 286 337
rect 288 335 290 337
rect 314 336 316 340
rect 325 336 327 340
rect 284 333 290 335
rect 274 331 280 333
rect 243 327 245 330
rect 257 327 259 330
rect 275 327 277 331
rect 175 309 177 314
rect 212 309 214 314
rect 33 295 90 297
rect 123 300 125 305
rect 133 297 135 305
rect 143 301 145 305
rect 157 301 159 305
rect 188 297 190 309
rect 288 319 290 333
rect 310 334 316 336
rect 310 332 312 334
rect 314 332 316 334
rect 310 330 316 332
rect 321 334 327 336
rect 335 337 337 340
rect 335 335 349 337
rect 321 332 323 334
rect 325 332 327 334
rect 321 330 327 332
rect 343 334 349 335
rect 343 332 345 334
rect 347 332 349 334
rect 312 327 314 330
rect 323 327 325 330
rect 333 327 335 331
rect 343 330 349 332
rect 355 336 357 342
rect 375 337 377 342
rect 388 339 390 342
rect 455 353 457 357
rect 445 341 447 345
rect 475 352 477 357
rect 488 349 490 361
rect 545 361 590 363
rect 545 356 547 361
rect 514 350 516 354
rect 525 351 527 356
rect 535 351 537 356
rect 384 337 390 339
rect 355 334 364 336
rect 355 332 360 334
rect 362 332 364 334
rect 355 330 364 332
rect 374 335 380 337
rect 374 333 376 335
rect 378 333 380 335
rect 384 335 386 337
rect 388 335 390 337
rect 414 336 416 340
rect 425 336 427 340
rect 384 333 390 335
rect 374 331 380 333
rect 343 327 345 330
rect 357 327 359 330
rect 375 327 377 331
rect 275 309 277 314
rect 312 309 314 314
rect 133 295 190 297
rect 223 300 225 305
rect 233 297 235 305
rect 243 301 245 305
rect 257 301 259 305
rect 288 297 290 309
rect 388 319 390 333
rect 410 334 416 336
rect 410 332 412 334
rect 414 332 416 334
rect 410 330 416 332
rect 421 334 427 336
rect 435 337 437 340
rect 435 335 449 337
rect 421 332 423 334
rect 425 332 427 334
rect 421 330 427 332
rect 443 334 449 335
rect 443 332 445 334
rect 447 332 449 334
rect 412 327 414 330
rect 423 327 425 330
rect 433 327 435 331
rect 443 330 449 332
rect 455 336 457 342
rect 475 337 477 342
rect 488 339 490 342
rect 555 353 557 357
rect 545 341 547 345
rect 575 352 577 357
rect 588 349 590 361
rect 645 361 690 363
rect 645 356 647 361
rect 614 350 616 354
rect 625 351 627 356
rect 635 351 637 356
rect 484 337 490 339
rect 455 334 464 336
rect 455 332 460 334
rect 462 332 464 334
rect 455 330 464 332
rect 474 335 480 337
rect 474 333 476 335
rect 478 333 480 335
rect 484 335 486 337
rect 488 335 490 337
rect 514 336 516 340
rect 525 336 527 340
rect 484 333 490 335
rect 474 331 480 333
rect 443 327 445 330
rect 457 327 459 330
rect 475 327 477 331
rect 375 309 377 314
rect 412 309 414 314
rect 233 295 290 297
rect 323 300 325 305
rect 333 297 335 305
rect 343 301 345 305
rect 357 301 359 305
rect 388 297 390 309
rect 488 319 490 333
rect 510 334 516 336
rect 510 332 512 334
rect 514 332 516 334
rect 510 330 516 332
rect 521 334 527 336
rect 535 337 537 340
rect 535 335 549 337
rect 521 332 523 334
rect 525 332 527 334
rect 521 330 527 332
rect 543 334 549 335
rect 543 332 545 334
rect 547 332 549 334
rect 512 327 514 330
rect 523 327 525 330
rect 533 327 535 331
rect 543 330 549 332
rect 555 336 557 342
rect 575 337 577 342
rect 588 339 590 342
rect 655 353 657 357
rect 645 341 647 345
rect 675 352 677 357
rect 688 349 690 361
rect 745 361 790 363
rect 745 356 747 361
rect 714 350 716 354
rect 725 351 727 356
rect 735 351 737 356
rect 584 337 590 339
rect 555 334 564 336
rect 555 332 560 334
rect 562 332 564 334
rect 555 330 564 332
rect 574 335 580 337
rect 574 333 576 335
rect 578 333 580 335
rect 584 335 586 337
rect 588 335 590 337
rect 614 336 616 340
rect 625 336 627 340
rect 584 333 590 335
rect 574 331 580 333
rect 543 327 545 330
rect 557 327 559 330
rect 575 327 577 331
rect 475 309 477 314
rect 512 309 514 314
rect 333 295 390 297
rect 423 300 425 305
rect 433 297 435 305
rect 443 301 445 305
rect 457 301 459 305
rect 488 297 490 309
rect 588 319 590 333
rect 610 334 616 336
rect 610 332 612 334
rect 614 332 616 334
rect 610 330 616 332
rect 621 334 627 336
rect 635 337 637 340
rect 635 335 649 337
rect 621 332 623 334
rect 625 332 627 334
rect 621 330 627 332
rect 643 334 649 335
rect 643 332 645 334
rect 647 332 649 334
rect 612 327 614 330
rect 623 327 625 330
rect 633 327 635 331
rect 643 330 649 332
rect 655 336 657 342
rect 675 337 677 342
rect 688 339 690 342
rect 755 353 757 357
rect 745 341 747 345
rect 775 352 777 357
rect 788 349 790 361
rect 684 337 690 339
rect 655 334 664 336
rect 655 332 660 334
rect 662 332 664 334
rect 655 330 664 332
rect 674 335 680 337
rect 674 333 676 335
rect 678 333 680 335
rect 684 335 686 337
rect 688 335 690 337
rect 714 336 716 340
rect 725 336 727 340
rect 684 333 690 335
rect 674 331 680 333
rect 643 327 645 330
rect 657 327 659 330
rect 675 327 677 331
rect 575 309 577 314
rect 612 309 614 314
rect 433 295 490 297
rect 523 300 525 305
rect 533 297 535 305
rect 543 301 545 305
rect 557 301 559 305
rect 588 297 590 309
rect 688 319 690 333
rect 710 334 716 336
rect 710 332 712 334
rect 714 332 716 334
rect 710 330 716 332
rect 721 334 727 336
rect 735 337 737 340
rect 735 335 749 337
rect 721 332 723 334
rect 725 332 727 334
rect 721 330 727 332
rect 743 334 749 335
rect 743 332 745 334
rect 747 332 749 334
rect 712 327 714 330
rect 723 327 725 330
rect 733 327 735 331
rect 743 330 749 332
rect 755 336 757 342
rect 775 337 777 342
rect 788 339 790 342
rect 784 337 790 339
rect 755 334 764 336
rect 755 332 760 334
rect 762 332 764 334
rect 755 330 764 332
rect 774 335 780 337
rect 774 333 776 335
rect 778 333 780 335
rect 784 335 786 337
rect 788 335 790 337
rect 784 333 790 335
rect 774 331 780 333
rect 743 327 745 330
rect 757 327 759 330
rect 775 327 777 331
rect 675 309 677 314
rect 712 309 714 314
rect 533 295 590 297
rect 623 300 625 305
rect 633 297 635 305
rect 643 301 645 305
rect 657 301 659 305
rect 688 297 690 309
rect 788 319 790 333
rect 775 309 777 314
rect 633 295 690 297
rect 723 300 725 305
rect 733 297 735 305
rect 743 301 745 305
rect 757 301 759 305
rect 788 297 790 309
rect 733 295 790 297
rect 12 289 69 291
rect 12 277 14 289
rect 43 281 45 285
rect 57 281 59 285
rect 67 281 69 289
rect 77 281 79 286
rect 112 289 169 291
rect 25 272 27 277
rect 12 253 14 267
rect 112 277 114 289
rect 143 281 145 285
rect 157 281 159 285
rect 167 281 169 289
rect 177 281 179 286
rect 212 289 269 291
rect 88 272 90 277
rect 125 272 127 277
rect 25 255 27 259
rect 43 256 45 259
rect 57 256 59 259
rect 22 253 28 255
rect 12 251 18 253
rect 12 249 14 251
rect 16 249 18 251
rect 22 251 24 253
rect 26 251 28 253
rect 22 249 28 251
rect 38 254 47 256
rect 38 252 40 254
rect 42 252 47 254
rect 38 250 47 252
rect 12 247 18 249
rect 12 244 14 247
rect 25 244 27 249
rect 45 244 47 250
rect 53 254 59 256
rect 67 255 69 259
rect 77 256 79 259
rect 88 256 90 259
rect 53 252 55 254
rect 57 252 59 254
rect 53 251 59 252
rect 75 254 81 256
rect 75 252 77 254
rect 79 252 81 254
rect 53 249 67 251
rect 65 246 67 249
rect 75 250 81 252
rect 86 254 92 256
rect 86 252 88 254
rect 90 252 92 254
rect 86 250 92 252
rect 112 253 114 267
rect 212 277 214 289
rect 243 281 245 285
rect 257 281 259 285
rect 267 281 269 289
rect 277 281 279 286
rect 312 289 369 291
rect 188 272 190 277
rect 225 272 227 277
rect 125 255 127 259
rect 143 256 145 259
rect 157 256 159 259
rect 122 253 128 255
rect 112 251 118 253
rect 75 246 77 250
rect 86 246 88 250
rect 112 249 114 251
rect 116 249 118 251
rect 122 251 124 253
rect 126 251 128 253
rect 122 249 128 251
rect 138 254 147 256
rect 138 252 140 254
rect 142 252 147 254
rect 138 250 147 252
rect 112 247 118 249
rect 12 225 14 237
rect 25 229 27 234
rect 55 241 57 245
rect 45 229 47 233
rect 112 244 114 247
rect 125 244 127 249
rect 145 244 147 250
rect 153 254 159 256
rect 167 255 169 259
rect 177 256 179 259
rect 188 256 190 259
rect 153 252 155 254
rect 157 252 159 254
rect 153 251 159 252
rect 175 254 181 256
rect 175 252 177 254
rect 179 252 181 254
rect 153 249 167 251
rect 165 246 167 249
rect 175 250 181 252
rect 186 254 192 256
rect 186 252 188 254
rect 190 252 192 254
rect 186 250 192 252
rect 212 253 214 267
rect 312 277 314 289
rect 343 281 345 285
rect 357 281 359 285
rect 367 281 369 289
rect 377 281 379 286
rect 414 289 471 291
rect 288 273 290 277
rect 325 272 327 277
rect 225 255 227 259
rect 243 256 245 259
rect 257 256 259 259
rect 222 253 228 255
rect 212 251 218 253
rect 175 246 177 250
rect 186 246 188 250
rect 212 249 214 251
rect 216 249 218 251
rect 222 251 224 253
rect 226 251 228 253
rect 222 249 228 251
rect 238 254 247 256
rect 238 252 240 254
rect 242 252 247 254
rect 238 250 247 252
rect 212 247 218 249
rect 65 230 67 235
rect 75 230 77 235
rect 86 232 88 236
rect 55 225 57 230
rect 12 223 57 225
rect 112 225 114 237
rect 125 229 127 234
rect 155 241 157 245
rect 145 229 147 233
rect 212 244 214 247
rect 225 244 227 249
rect 245 244 247 250
rect 253 254 259 256
rect 267 255 269 259
rect 277 256 279 259
rect 288 256 290 259
rect 253 252 255 254
rect 257 252 259 254
rect 253 251 259 252
rect 275 254 281 256
rect 275 252 277 254
rect 279 252 281 254
rect 253 249 267 251
rect 265 246 267 249
rect 275 250 281 252
rect 286 254 292 256
rect 286 252 288 254
rect 290 252 292 254
rect 286 250 292 252
rect 312 253 314 267
rect 414 277 416 289
rect 445 281 447 285
rect 459 281 461 285
rect 469 281 471 289
rect 479 281 481 286
rect 514 289 571 291
rect 388 272 390 277
rect 427 272 429 277
rect 325 255 327 259
rect 343 256 345 259
rect 357 256 359 259
rect 322 253 328 255
rect 312 251 318 253
rect 275 246 277 250
rect 286 246 288 250
rect 312 249 314 251
rect 316 249 318 251
rect 322 251 324 253
rect 326 251 328 253
rect 322 249 328 251
rect 338 254 347 256
rect 338 252 340 254
rect 342 252 347 254
rect 338 250 347 252
rect 312 247 318 249
rect 165 230 167 235
rect 175 230 177 235
rect 186 232 188 236
rect 155 225 157 230
rect 112 223 157 225
rect 212 225 214 237
rect 225 229 227 234
rect 255 241 257 245
rect 245 229 247 233
rect 312 244 314 247
rect 325 244 327 249
rect 345 244 347 250
rect 353 254 359 256
rect 367 255 369 259
rect 377 256 379 259
rect 388 256 390 259
rect 353 252 355 254
rect 357 252 359 254
rect 353 251 359 252
rect 375 254 381 256
rect 375 252 377 254
rect 379 252 381 254
rect 353 249 367 251
rect 365 246 367 249
rect 375 250 381 252
rect 386 254 392 256
rect 386 252 388 254
rect 390 252 392 254
rect 386 250 392 252
rect 414 253 416 267
rect 514 277 516 289
rect 545 281 547 285
rect 559 281 561 285
rect 569 281 571 289
rect 579 281 581 286
rect 614 289 671 291
rect 490 273 492 277
rect 527 272 529 277
rect 427 255 429 259
rect 445 256 447 259
rect 459 256 461 259
rect 424 253 430 255
rect 414 251 420 253
rect 375 246 377 250
rect 386 246 388 250
rect 414 249 416 251
rect 418 249 420 251
rect 424 251 426 253
rect 428 251 430 253
rect 424 249 430 251
rect 440 254 449 256
rect 440 252 442 254
rect 444 252 449 254
rect 440 250 449 252
rect 414 247 420 249
rect 265 230 267 235
rect 275 230 277 235
rect 286 232 288 236
rect 255 225 257 230
rect 212 223 257 225
rect 312 225 314 237
rect 325 229 327 234
rect 355 241 357 245
rect 345 229 347 233
rect 414 244 416 247
rect 427 244 429 249
rect 447 244 449 250
rect 455 254 461 256
rect 469 255 471 259
rect 479 256 481 259
rect 490 256 492 260
rect 455 252 457 254
rect 459 252 461 254
rect 455 251 461 252
rect 477 254 483 256
rect 477 252 479 254
rect 481 252 483 254
rect 455 249 469 251
rect 467 246 469 249
rect 477 250 483 252
rect 488 254 494 256
rect 488 252 490 254
rect 492 252 494 254
rect 488 250 494 252
rect 514 253 516 267
rect 614 277 616 289
rect 645 281 647 285
rect 659 281 661 285
rect 669 281 671 289
rect 679 281 681 286
rect 714 289 771 291
rect 590 272 592 277
rect 627 272 629 277
rect 527 255 529 259
rect 545 256 547 259
rect 559 256 561 259
rect 524 253 530 255
rect 514 251 520 253
rect 477 246 479 250
rect 488 246 490 250
rect 514 249 516 251
rect 518 249 520 251
rect 524 251 526 253
rect 528 251 530 253
rect 524 249 530 251
rect 540 254 549 256
rect 540 252 542 254
rect 544 252 549 254
rect 540 250 549 252
rect 514 247 520 249
rect 365 230 367 235
rect 375 230 377 235
rect 386 232 388 236
rect 355 225 357 230
rect 312 223 357 225
rect 414 225 416 237
rect 427 229 429 234
rect 457 241 459 245
rect 447 229 449 233
rect 514 244 516 247
rect 527 244 529 249
rect 547 244 549 250
rect 555 254 561 256
rect 569 255 571 259
rect 579 256 581 259
rect 590 256 592 259
rect 555 252 557 254
rect 559 252 561 254
rect 555 251 561 252
rect 577 254 583 256
rect 577 252 579 254
rect 581 252 583 254
rect 555 249 569 251
rect 567 246 569 249
rect 577 250 583 252
rect 588 254 594 256
rect 588 252 590 254
rect 592 252 594 254
rect 588 250 594 252
rect 614 253 616 267
rect 714 277 716 289
rect 745 281 747 285
rect 759 281 761 285
rect 769 281 771 289
rect 779 281 781 286
rect 690 273 692 277
rect 727 272 729 277
rect 627 255 629 259
rect 645 256 647 259
rect 659 256 661 259
rect 624 253 630 255
rect 614 251 620 253
rect 577 246 579 250
rect 588 246 590 250
rect 614 249 616 251
rect 618 249 620 251
rect 624 251 626 253
rect 628 251 630 253
rect 624 249 630 251
rect 640 254 649 256
rect 640 252 642 254
rect 644 252 649 254
rect 640 250 649 252
rect 614 247 620 249
rect 467 230 469 235
rect 477 230 479 235
rect 488 232 490 236
rect 457 225 459 230
rect 414 223 459 225
rect 514 225 516 237
rect 527 229 529 234
rect 557 241 559 245
rect 547 229 549 233
rect 614 244 616 247
rect 627 244 629 249
rect 647 244 649 250
rect 655 254 661 256
rect 669 255 671 259
rect 679 256 681 259
rect 690 256 692 260
rect 655 252 657 254
rect 659 252 661 254
rect 655 251 661 252
rect 677 254 683 256
rect 677 252 679 254
rect 681 252 683 254
rect 655 249 669 251
rect 667 246 669 249
rect 677 250 683 252
rect 688 254 694 256
rect 688 252 690 254
rect 692 252 694 254
rect 688 250 694 252
rect 714 253 716 267
rect 790 272 792 277
rect 727 255 729 259
rect 745 256 747 259
rect 759 256 761 259
rect 724 253 730 255
rect 714 251 720 253
rect 677 246 679 250
rect 688 246 690 250
rect 714 249 716 251
rect 718 249 720 251
rect 724 251 726 253
rect 728 251 730 253
rect 724 249 730 251
rect 740 254 749 256
rect 740 252 742 254
rect 744 252 749 254
rect 740 250 749 252
rect 714 247 720 249
rect 567 230 569 235
rect 577 230 579 235
rect 588 232 590 236
rect 557 225 559 230
rect 514 223 559 225
rect 614 225 616 237
rect 627 229 629 234
rect 657 241 659 245
rect 647 229 649 233
rect 714 244 716 247
rect 727 244 729 249
rect 747 244 749 250
rect 755 254 761 256
rect 769 255 771 259
rect 779 256 781 259
rect 790 256 792 259
rect 755 252 757 254
rect 759 252 761 254
rect 755 251 761 252
rect 777 254 783 256
rect 777 252 779 254
rect 781 252 783 254
rect 755 249 769 251
rect 767 246 769 249
rect 777 250 783 252
rect 788 254 794 256
rect 788 252 790 254
rect 792 252 794 254
rect 788 250 794 252
rect 777 246 779 250
rect 788 246 790 250
rect 667 230 669 235
rect 677 230 679 235
rect 688 232 690 236
rect 657 225 659 230
rect 614 223 659 225
rect 714 225 716 237
rect 727 229 729 234
rect 757 241 759 245
rect 747 229 749 233
rect 767 230 769 235
rect 777 230 779 235
rect 788 232 790 236
rect 757 225 759 230
rect 714 223 759 225
rect 12 217 57 219
rect 12 205 14 217
rect 25 208 27 213
rect 45 209 47 213
rect 55 212 57 217
rect 112 217 157 219
rect 65 207 67 212
rect 75 207 77 212
rect 12 195 14 198
rect 12 193 18 195
rect 25 193 27 198
rect 12 191 14 193
rect 16 191 18 193
rect 12 189 18 191
rect 22 191 28 193
rect 45 192 47 198
rect 55 197 57 201
rect 86 206 88 210
rect 112 205 114 217
rect 125 208 127 213
rect 145 209 147 213
rect 155 212 157 217
rect 212 217 257 219
rect 165 207 167 212
rect 175 207 177 212
rect 65 193 67 196
rect 22 189 24 191
rect 26 189 28 191
rect 12 175 14 189
rect 22 187 28 189
rect 38 190 47 192
rect 38 188 40 190
rect 42 188 47 190
rect 25 183 27 187
rect 38 186 47 188
rect 53 191 67 193
rect 75 192 77 196
rect 86 192 88 196
rect 112 195 114 198
rect 112 193 118 195
rect 125 194 127 198
rect 53 190 59 191
rect 53 188 55 190
rect 57 188 59 190
rect 53 186 59 188
rect 75 190 81 192
rect 75 188 77 190
rect 79 188 81 190
rect 43 183 45 186
rect 57 183 59 186
rect 67 183 69 187
rect 75 186 81 188
rect 86 190 92 192
rect 86 188 88 190
rect 90 188 92 190
rect 86 186 92 188
rect 112 191 114 193
rect 116 191 118 193
rect 112 189 118 191
rect 122 192 128 194
rect 145 192 147 198
rect 155 197 157 201
rect 186 206 188 210
rect 212 205 214 217
rect 225 208 227 213
rect 245 209 247 213
rect 255 212 257 217
rect 312 217 357 219
rect 265 207 267 212
rect 275 207 277 212
rect 165 193 167 196
rect 122 190 124 192
rect 126 190 128 192
rect 77 183 79 186
rect 88 183 90 186
rect 25 165 27 170
rect 12 153 14 165
rect 112 175 114 189
rect 122 188 128 190
rect 138 190 147 192
rect 138 188 140 190
rect 142 188 147 190
rect 125 183 127 188
rect 138 186 147 188
rect 153 191 167 193
rect 175 192 177 196
rect 186 192 188 196
rect 212 195 214 198
rect 212 193 218 195
rect 225 193 227 198
rect 153 190 159 191
rect 153 188 155 190
rect 157 188 159 190
rect 153 186 159 188
rect 175 190 181 192
rect 175 188 177 190
rect 179 188 181 190
rect 143 183 145 186
rect 157 183 159 186
rect 167 183 169 187
rect 175 186 181 188
rect 186 190 192 192
rect 186 188 188 190
rect 190 188 192 190
rect 186 186 192 188
rect 212 191 214 193
rect 216 191 218 193
rect 212 189 218 191
rect 222 191 228 193
rect 245 192 247 198
rect 255 197 257 201
rect 286 206 288 210
rect 312 205 314 217
rect 325 208 327 213
rect 345 209 347 213
rect 355 212 357 217
rect 414 217 459 219
rect 365 207 367 212
rect 375 207 377 212
rect 265 193 267 196
rect 222 189 224 191
rect 226 189 228 191
rect 177 183 179 186
rect 188 183 190 186
rect 88 165 90 170
rect 125 165 127 170
rect 43 157 45 161
rect 57 157 59 161
rect 67 153 69 161
rect 77 156 79 161
rect 12 151 69 153
rect 112 153 114 165
rect 212 175 214 189
rect 222 187 228 189
rect 238 190 247 192
rect 238 188 240 190
rect 242 188 247 190
rect 225 183 227 187
rect 238 186 247 188
rect 253 191 267 193
rect 275 192 277 196
rect 286 192 288 196
rect 312 195 314 198
rect 312 193 318 195
rect 325 194 327 198
rect 253 190 259 191
rect 253 188 255 190
rect 257 188 259 190
rect 253 186 259 188
rect 275 190 281 192
rect 275 188 277 190
rect 279 188 281 190
rect 243 183 245 186
rect 257 183 259 186
rect 267 183 269 187
rect 275 186 281 188
rect 286 190 292 192
rect 286 188 288 190
rect 290 188 292 190
rect 286 186 292 188
rect 312 191 314 193
rect 316 191 318 193
rect 312 189 318 191
rect 322 192 328 194
rect 345 192 347 198
rect 355 197 357 201
rect 386 206 388 210
rect 414 205 416 217
rect 427 208 429 213
rect 447 209 449 213
rect 457 212 459 217
rect 514 217 559 219
rect 467 207 469 212
rect 477 207 479 212
rect 365 193 367 196
rect 322 190 324 192
rect 326 190 328 192
rect 277 183 279 186
rect 288 183 290 186
rect 188 165 190 170
rect 225 165 227 170
rect 143 157 145 161
rect 157 157 159 161
rect 167 153 169 161
rect 177 156 179 161
rect 112 151 169 153
rect 212 153 214 165
rect 312 175 314 189
rect 322 188 328 190
rect 338 190 347 192
rect 338 188 340 190
rect 342 188 347 190
rect 325 183 327 188
rect 338 186 347 188
rect 353 191 367 193
rect 375 192 377 196
rect 386 192 388 196
rect 414 195 416 198
rect 414 193 420 195
rect 427 193 429 198
rect 353 190 359 191
rect 353 188 355 190
rect 357 188 359 190
rect 353 186 359 188
rect 375 190 381 192
rect 375 188 377 190
rect 379 188 381 190
rect 343 183 345 186
rect 357 183 359 186
rect 367 183 369 187
rect 375 186 381 188
rect 385 190 392 192
rect 385 188 387 190
rect 389 188 392 190
rect 385 186 392 188
rect 414 191 416 193
rect 418 191 420 193
rect 414 189 420 191
rect 424 191 430 193
rect 447 192 449 198
rect 457 197 459 201
rect 488 206 490 210
rect 514 205 516 217
rect 527 208 529 213
rect 547 209 549 213
rect 557 212 559 217
rect 614 217 659 219
rect 567 207 569 212
rect 577 207 579 212
rect 467 193 469 196
rect 424 189 426 191
rect 428 189 430 191
rect 377 183 379 186
rect 388 183 390 186
rect 288 165 290 170
rect 325 165 327 170
rect 243 157 245 161
rect 257 157 259 161
rect 267 153 269 161
rect 277 156 279 161
rect 212 151 269 153
rect 312 153 314 165
rect 414 175 416 189
rect 424 187 430 189
rect 440 190 449 192
rect 440 188 442 190
rect 444 188 449 190
rect 427 183 429 187
rect 440 186 449 188
rect 455 191 469 193
rect 477 192 479 196
rect 488 192 490 196
rect 514 195 516 198
rect 514 193 520 195
rect 527 194 529 198
rect 455 190 461 191
rect 455 188 457 190
rect 459 188 461 190
rect 455 186 461 188
rect 477 190 483 192
rect 477 188 479 190
rect 481 188 483 190
rect 445 183 447 186
rect 459 183 461 186
rect 469 183 471 187
rect 477 186 483 188
rect 488 190 494 192
rect 488 188 490 190
rect 492 188 494 190
rect 488 186 494 188
rect 514 191 516 193
rect 518 191 520 193
rect 514 189 520 191
rect 524 192 530 194
rect 547 192 549 198
rect 557 197 559 201
rect 588 206 590 210
rect 614 205 616 217
rect 627 208 629 213
rect 647 209 649 213
rect 657 212 659 217
rect 714 217 759 219
rect 667 207 669 212
rect 677 207 679 212
rect 567 193 569 196
rect 524 190 526 192
rect 528 190 530 192
rect 479 183 481 186
rect 490 183 492 186
rect 388 165 390 170
rect 427 165 429 170
rect 343 157 345 161
rect 357 157 359 161
rect 367 153 369 161
rect 377 156 379 161
rect 312 151 369 153
rect 414 153 416 165
rect 514 175 516 189
rect 524 188 530 190
rect 540 190 549 192
rect 540 188 542 190
rect 544 188 549 190
rect 527 183 529 188
rect 540 186 549 188
rect 555 191 569 193
rect 577 192 579 196
rect 588 192 590 196
rect 614 195 616 198
rect 614 193 620 195
rect 627 193 629 198
rect 555 190 561 191
rect 555 188 557 190
rect 559 188 561 190
rect 555 186 561 188
rect 577 190 583 192
rect 577 188 579 190
rect 581 188 583 190
rect 545 183 547 186
rect 559 183 561 186
rect 569 183 571 187
rect 577 186 583 188
rect 588 190 594 192
rect 588 188 590 190
rect 592 188 594 190
rect 588 186 594 188
rect 614 191 616 193
rect 618 191 620 193
rect 614 189 620 191
rect 624 191 630 193
rect 647 192 649 198
rect 657 197 659 201
rect 688 206 690 210
rect 714 205 716 217
rect 727 208 729 213
rect 747 209 749 213
rect 757 212 759 217
rect 767 207 769 212
rect 777 207 779 212
rect 667 193 669 196
rect 624 189 626 191
rect 628 189 630 191
rect 579 183 581 186
rect 590 183 592 186
rect 490 165 492 170
rect 527 165 529 170
rect 445 157 447 161
rect 459 157 461 161
rect 469 153 471 161
rect 479 156 481 161
rect 414 151 471 153
rect 514 153 516 165
rect 614 175 616 189
rect 624 187 630 189
rect 640 190 649 192
rect 640 188 642 190
rect 644 188 649 190
rect 627 183 629 187
rect 640 186 649 188
rect 655 191 669 193
rect 677 192 679 196
rect 688 192 690 196
rect 714 195 716 198
rect 714 193 720 195
rect 727 194 729 198
rect 655 190 661 191
rect 655 188 657 190
rect 659 188 661 190
rect 655 186 661 188
rect 677 190 683 192
rect 677 188 679 190
rect 681 188 683 190
rect 645 183 647 186
rect 659 183 661 186
rect 669 183 671 187
rect 677 186 683 188
rect 688 190 694 192
rect 688 188 690 190
rect 692 188 694 190
rect 688 186 694 188
rect 714 191 716 193
rect 718 191 720 193
rect 714 189 720 191
rect 724 192 730 194
rect 747 192 749 198
rect 757 197 759 201
rect 788 206 790 210
rect 767 193 769 196
rect 724 190 726 192
rect 728 190 730 192
rect 679 183 681 186
rect 690 183 692 186
rect 590 165 592 170
rect 627 165 629 170
rect 545 157 547 161
rect 559 157 561 161
rect 569 153 571 161
rect 579 156 581 161
rect 514 151 571 153
rect 614 153 616 165
rect 714 175 716 189
rect 724 188 730 190
rect 740 190 749 192
rect 740 188 742 190
rect 744 188 749 190
rect 727 183 729 188
rect 740 186 749 188
rect 755 191 769 193
rect 777 192 779 196
rect 788 192 790 196
rect 755 190 761 191
rect 755 188 757 190
rect 759 188 761 190
rect 755 186 761 188
rect 777 190 783 192
rect 777 188 779 190
rect 781 188 783 190
rect 745 183 747 186
rect 759 183 761 186
rect 769 183 771 187
rect 777 186 783 188
rect 788 190 794 192
rect 788 188 790 190
rect 792 188 794 190
rect 788 186 794 188
rect 779 183 781 186
rect 790 183 792 186
rect 690 165 692 170
rect 727 165 729 170
rect 645 157 647 161
rect 659 157 661 161
rect 669 153 671 161
rect 679 156 681 161
rect 614 151 671 153
rect 714 153 716 165
rect 790 165 792 170
rect 745 157 747 161
rect 759 157 761 161
rect 769 153 771 161
rect 779 156 781 161
rect 714 151 771 153
rect 12 145 69 147
rect 12 133 14 145
rect 43 137 45 141
rect 57 137 59 141
rect 67 137 69 145
rect 77 137 79 142
rect 112 145 169 147
rect 25 128 27 133
rect 12 109 14 123
rect 112 133 114 145
rect 143 137 145 141
rect 157 137 159 141
rect 167 137 169 145
rect 177 137 179 142
rect 212 145 269 147
rect 88 128 90 133
rect 125 128 127 133
rect 25 111 27 115
rect 43 112 45 115
rect 57 112 59 115
rect 22 109 28 111
rect 12 107 18 109
rect 12 105 14 107
rect 16 105 18 107
rect 22 107 24 109
rect 26 107 28 109
rect 22 105 28 107
rect 38 110 47 112
rect 38 108 40 110
rect 42 108 47 110
rect 38 106 47 108
rect 12 103 18 105
rect 12 100 14 103
rect 25 100 27 105
rect 45 100 47 106
rect 53 110 59 112
rect 67 111 69 115
rect 77 112 79 115
rect 88 112 90 115
rect 53 108 55 110
rect 57 108 59 110
rect 53 107 59 108
rect 75 110 81 112
rect 75 108 77 110
rect 79 108 81 110
rect 53 105 67 107
rect 65 102 67 105
rect 75 106 81 108
rect 86 110 92 112
rect 86 108 88 110
rect 90 108 92 110
rect 86 106 92 108
rect 112 109 114 123
rect 212 133 214 145
rect 243 137 245 141
rect 257 137 259 141
rect 267 137 269 145
rect 277 137 279 142
rect 312 145 369 147
rect 188 128 190 133
rect 225 128 227 133
rect 125 111 127 115
rect 143 112 145 115
rect 157 112 159 115
rect 123 109 129 111
rect 112 107 118 109
rect 75 102 77 106
rect 86 102 88 106
rect 112 105 114 107
rect 116 105 118 107
rect 123 107 125 109
rect 127 107 129 109
rect 123 105 129 107
rect 138 110 147 112
rect 138 108 140 110
rect 142 108 147 110
rect 138 106 147 108
rect 112 103 118 105
rect 12 81 14 93
rect 25 85 27 90
rect 55 97 57 101
rect 45 85 47 89
rect 112 100 114 103
rect 125 100 127 105
rect 145 100 147 106
rect 153 110 159 112
rect 167 111 169 115
rect 177 112 179 115
rect 188 112 190 115
rect 153 108 155 110
rect 157 108 159 110
rect 153 107 159 108
rect 175 110 181 112
rect 175 108 177 110
rect 179 108 181 110
rect 153 105 167 107
rect 165 102 167 105
rect 175 106 181 108
rect 186 110 192 112
rect 186 108 188 110
rect 190 108 192 110
rect 186 106 192 108
rect 212 109 214 123
rect 312 133 314 145
rect 343 137 345 141
rect 357 137 359 141
rect 367 137 369 145
rect 377 137 379 142
rect 414 145 471 147
rect 288 128 290 133
rect 325 128 327 133
rect 225 111 227 115
rect 243 112 245 115
rect 257 112 259 115
rect 222 109 228 111
rect 212 107 218 109
rect 175 102 177 106
rect 186 102 188 106
rect 212 105 214 107
rect 216 105 218 107
rect 222 107 224 109
rect 226 107 228 109
rect 222 105 228 107
rect 238 110 247 112
rect 238 108 240 110
rect 242 108 247 110
rect 238 106 247 108
rect 212 103 218 105
rect 65 86 67 91
rect 75 86 77 91
rect 86 88 88 92
rect 55 81 57 86
rect 12 79 57 81
rect 112 81 114 93
rect 125 85 127 90
rect 155 97 157 101
rect 145 85 147 89
rect 212 100 214 103
rect 225 100 227 105
rect 245 100 247 106
rect 253 110 259 112
rect 267 111 269 115
rect 277 112 279 115
rect 288 112 290 115
rect 253 108 255 110
rect 257 108 259 110
rect 253 107 259 108
rect 275 110 281 112
rect 275 108 277 110
rect 279 108 281 110
rect 253 105 267 107
rect 265 102 267 105
rect 275 106 281 108
rect 286 110 292 112
rect 286 108 288 110
rect 290 108 292 110
rect 286 106 292 108
rect 312 109 314 123
rect 414 133 416 145
rect 445 137 447 141
rect 459 137 461 141
rect 469 137 471 145
rect 479 137 481 142
rect 514 145 571 147
rect 388 128 390 133
rect 427 128 429 133
rect 325 111 327 115
rect 343 112 345 115
rect 357 112 359 115
rect 322 109 328 111
rect 312 107 318 109
rect 275 102 277 106
rect 286 102 288 106
rect 312 105 314 107
rect 316 105 318 107
rect 322 107 324 109
rect 326 107 328 109
rect 322 105 328 107
rect 338 110 347 112
rect 338 108 340 110
rect 342 108 347 110
rect 338 106 347 108
rect 312 103 318 105
rect 165 86 167 91
rect 175 86 177 91
rect 186 88 188 92
rect 155 81 157 86
rect 112 79 157 81
rect 212 81 214 93
rect 225 85 227 90
rect 255 97 257 101
rect 245 85 247 89
rect 312 100 314 103
rect 325 100 327 105
rect 345 100 347 106
rect 353 110 359 112
rect 367 111 369 115
rect 377 112 379 115
rect 388 112 390 115
rect 353 108 355 110
rect 357 108 359 110
rect 353 107 359 108
rect 375 110 381 112
rect 375 108 377 110
rect 379 108 381 110
rect 353 105 367 107
rect 365 102 367 105
rect 375 106 381 108
rect 386 110 392 112
rect 386 108 388 110
rect 390 108 392 110
rect 386 106 392 108
rect 414 109 416 123
rect 514 133 516 145
rect 545 137 547 141
rect 559 137 561 141
rect 569 137 571 145
rect 579 137 581 142
rect 614 145 671 147
rect 490 128 492 133
rect 527 128 529 133
rect 427 111 429 115
rect 445 112 447 115
rect 459 112 461 115
rect 424 109 430 111
rect 414 107 420 109
rect 375 102 377 106
rect 386 102 388 106
rect 414 105 416 107
rect 418 105 420 107
rect 424 107 426 109
rect 428 107 430 109
rect 424 105 430 107
rect 440 110 449 112
rect 440 108 442 110
rect 444 108 449 110
rect 440 106 449 108
rect 414 103 420 105
rect 265 86 267 91
rect 275 86 277 91
rect 286 88 288 92
rect 255 81 257 86
rect 212 79 257 81
rect 312 81 314 93
rect 325 85 327 90
rect 355 97 357 101
rect 345 85 347 89
rect 414 100 416 103
rect 427 100 429 105
rect 447 100 449 106
rect 455 110 461 112
rect 469 111 471 115
rect 479 112 481 115
rect 490 112 492 115
rect 455 108 457 110
rect 459 108 461 110
rect 455 107 461 108
rect 477 110 483 112
rect 477 108 479 110
rect 481 108 483 110
rect 455 105 469 107
rect 467 102 469 105
rect 477 106 483 108
rect 488 110 494 112
rect 488 108 490 110
rect 492 108 494 110
rect 488 106 494 108
rect 514 109 516 123
rect 614 133 616 145
rect 645 137 647 141
rect 659 137 661 141
rect 669 137 671 145
rect 679 137 681 142
rect 714 145 771 147
rect 590 128 592 133
rect 627 128 629 133
rect 527 111 529 115
rect 545 112 547 115
rect 559 112 561 115
rect 524 109 530 111
rect 514 107 520 109
rect 477 102 479 106
rect 488 102 490 106
rect 514 105 516 107
rect 518 105 520 107
rect 524 107 526 109
rect 528 107 530 109
rect 524 105 530 107
rect 540 110 549 112
rect 540 108 542 110
rect 544 108 549 110
rect 540 106 549 108
rect 514 103 520 105
rect 365 86 367 91
rect 375 86 377 91
rect 386 88 388 92
rect 355 81 357 86
rect 312 79 357 81
rect 414 81 416 93
rect 427 85 429 90
rect 457 97 459 101
rect 447 85 449 89
rect 514 100 516 103
rect 527 100 529 105
rect 547 100 549 106
rect 555 110 561 112
rect 569 111 571 115
rect 579 112 581 115
rect 590 112 592 115
rect 555 108 557 110
rect 559 108 561 110
rect 555 107 561 108
rect 577 110 583 112
rect 577 108 579 110
rect 581 108 583 110
rect 555 105 569 107
rect 567 102 569 105
rect 577 106 583 108
rect 588 110 594 112
rect 588 108 590 110
rect 592 108 594 110
rect 588 106 594 108
rect 614 109 616 123
rect 714 133 716 145
rect 745 137 747 141
rect 759 137 761 141
rect 769 137 771 145
rect 779 137 781 142
rect 690 128 692 133
rect 727 128 729 133
rect 627 111 629 115
rect 645 112 647 115
rect 659 112 661 115
rect 624 109 630 111
rect 614 107 620 109
rect 577 102 579 106
rect 588 102 590 106
rect 614 105 616 107
rect 618 105 620 107
rect 624 107 626 109
rect 628 107 630 109
rect 624 105 630 107
rect 640 110 649 112
rect 640 108 642 110
rect 644 108 649 110
rect 640 106 649 108
rect 614 103 620 105
rect 467 86 469 91
rect 477 86 479 91
rect 488 88 490 92
rect 457 81 459 86
rect 414 79 459 81
rect 514 81 516 93
rect 527 85 529 90
rect 557 97 559 101
rect 547 85 549 89
rect 614 100 616 103
rect 627 100 629 105
rect 647 100 649 106
rect 655 110 661 112
rect 669 111 671 115
rect 679 112 681 115
rect 690 112 692 115
rect 655 108 657 110
rect 659 108 661 110
rect 655 107 661 108
rect 677 110 683 112
rect 677 108 679 110
rect 681 108 683 110
rect 655 105 669 107
rect 667 102 669 105
rect 677 106 683 108
rect 688 110 694 112
rect 688 108 690 110
rect 692 108 694 110
rect 688 106 694 108
rect 714 109 716 123
rect 790 128 792 133
rect 727 111 729 115
rect 745 112 747 115
rect 759 112 761 115
rect 724 109 730 111
rect 714 107 720 109
rect 677 102 679 106
rect 688 102 690 106
rect 714 105 716 107
rect 718 105 720 107
rect 724 107 726 109
rect 728 107 730 109
rect 724 105 730 107
rect 740 110 749 112
rect 740 108 742 110
rect 744 108 749 110
rect 740 106 749 108
rect 714 103 720 105
rect 567 86 569 91
rect 577 86 579 91
rect 588 88 590 92
rect 557 81 559 86
rect 514 79 559 81
rect 614 81 616 93
rect 627 85 629 90
rect 657 97 659 101
rect 647 85 649 89
rect 714 100 716 103
rect 727 100 729 105
rect 747 100 749 106
rect 755 110 761 112
rect 769 111 771 115
rect 779 112 781 115
rect 790 112 792 115
rect 755 108 757 110
rect 759 108 761 110
rect 755 107 761 108
rect 777 110 783 112
rect 777 108 779 110
rect 781 108 783 110
rect 755 105 769 107
rect 767 102 769 105
rect 777 106 783 108
rect 788 110 794 112
rect 788 108 790 110
rect 792 108 794 110
rect 788 106 794 108
rect 777 102 779 106
rect 788 102 790 106
rect 667 86 669 91
rect 677 86 679 91
rect 688 88 690 92
rect 657 81 659 86
rect 614 79 659 81
rect 714 81 716 93
rect 727 85 729 90
rect 757 97 759 101
rect 747 85 749 89
rect 767 86 769 91
rect 777 86 779 91
rect 788 88 790 92
rect 757 81 759 86
rect 714 79 759 81
rect 45 73 90 75
rect 45 68 47 73
rect 14 62 16 66
rect 25 63 27 68
rect 35 63 37 68
rect 55 65 57 69
rect 45 53 47 57
rect 75 64 77 69
rect 88 61 90 73
rect 145 73 190 75
rect 145 68 147 73
rect 114 62 116 66
rect 125 63 127 68
rect 135 63 137 68
rect 14 48 16 52
rect 25 48 27 52
rect 10 46 16 48
rect 10 44 12 46
rect 14 44 16 46
rect 10 42 16 44
rect 21 46 27 48
rect 35 49 37 52
rect 35 47 49 49
rect 21 44 23 46
rect 25 44 27 46
rect 21 42 27 44
rect 43 46 49 47
rect 43 44 45 46
rect 47 44 49 46
rect 12 39 14 42
rect 23 39 25 42
rect 33 39 35 43
rect 43 42 49 44
rect 55 48 57 54
rect 75 49 77 54
rect 88 51 90 54
rect 155 65 157 69
rect 145 53 147 57
rect 175 64 177 69
rect 188 61 190 73
rect 245 73 290 75
rect 245 68 247 73
rect 214 62 216 66
rect 225 63 227 68
rect 235 63 237 68
rect 84 49 90 51
rect 55 46 64 48
rect 55 44 60 46
rect 62 44 64 46
rect 55 42 64 44
rect 74 47 80 49
rect 74 45 76 47
rect 78 45 80 47
rect 84 47 86 49
rect 88 47 90 49
rect 114 48 116 52
rect 125 48 127 52
rect 84 45 90 47
rect 74 43 80 45
rect 43 39 45 42
rect 57 39 59 42
rect 75 39 77 43
rect 12 21 14 26
rect 88 31 90 45
rect 110 46 116 48
rect 110 44 112 46
rect 114 44 116 46
rect 110 42 116 44
rect 121 46 127 48
rect 135 49 137 52
rect 135 47 149 49
rect 121 44 123 46
rect 125 44 127 46
rect 121 42 127 44
rect 143 46 149 47
rect 143 44 145 46
rect 147 44 149 46
rect 112 39 114 42
rect 123 39 125 42
rect 133 39 135 43
rect 143 42 149 44
rect 155 48 157 54
rect 175 49 177 54
rect 188 51 190 54
rect 255 65 257 69
rect 245 53 247 57
rect 275 64 277 69
rect 288 61 290 73
rect 345 73 390 75
rect 345 68 347 73
rect 314 62 316 66
rect 325 63 327 68
rect 335 63 337 68
rect 184 49 190 51
rect 155 46 164 48
rect 155 44 160 46
rect 162 44 164 46
rect 155 42 164 44
rect 174 47 180 49
rect 174 45 176 47
rect 178 45 180 47
rect 184 47 186 49
rect 188 47 190 49
rect 214 48 216 52
rect 225 48 227 52
rect 184 45 190 47
rect 174 43 180 45
rect 143 39 145 42
rect 157 39 159 42
rect 175 39 177 43
rect 75 21 77 26
rect 112 21 114 26
rect 23 12 25 17
rect 33 9 35 17
rect 43 13 45 17
rect 57 13 59 17
rect 88 9 90 21
rect 188 31 190 45
rect 210 46 216 48
rect 210 44 212 46
rect 214 44 216 46
rect 210 42 216 44
rect 221 46 227 48
rect 235 49 237 52
rect 235 47 249 49
rect 221 44 223 46
rect 225 44 227 46
rect 221 42 227 44
rect 243 46 249 47
rect 243 44 245 46
rect 247 44 249 46
rect 212 39 214 42
rect 223 39 225 42
rect 233 39 235 43
rect 243 42 249 44
rect 255 48 257 54
rect 275 49 277 54
rect 288 51 290 54
rect 355 65 357 69
rect 345 53 347 57
rect 375 64 377 69
rect 388 61 390 73
rect 445 73 490 75
rect 445 68 447 73
rect 414 62 416 66
rect 425 63 427 68
rect 435 63 437 68
rect 284 49 290 51
rect 255 46 264 48
rect 255 44 260 46
rect 262 44 264 46
rect 255 42 264 44
rect 274 47 280 49
rect 274 45 276 47
rect 278 45 280 47
rect 284 47 286 49
rect 288 47 290 49
rect 314 48 316 52
rect 325 48 327 52
rect 284 45 290 47
rect 274 43 280 45
rect 243 39 245 42
rect 257 39 259 42
rect 275 39 277 43
rect 175 21 177 26
rect 212 21 214 26
rect 33 7 90 9
rect 123 12 125 17
rect 133 9 135 17
rect 143 13 145 17
rect 157 13 159 17
rect 188 9 190 21
rect 288 31 290 45
rect 310 46 316 48
rect 310 44 312 46
rect 314 44 316 46
rect 310 42 316 44
rect 321 46 327 48
rect 335 49 337 52
rect 335 47 349 49
rect 321 44 323 46
rect 325 44 327 46
rect 321 42 327 44
rect 343 46 349 47
rect 343 44 345 46
rect 347 44 349 46
rect 312 39 314 42
rect 323 39 325 42
rect 333 39 335 43
rect 343 42 349 44
rect 355 48 357 54
rect 375 49 377 54
rect 388 51 390 54
rect 455 65 457 69
rect 445 53 447 57
rect 475 64 477 69
rect 488 61 490 73
rect 545 73 590 75
rect 545 68 547 73
rect 514 62 516 66
rect 525 63 527 68
rect 535 63 537 68
rect 384 49 390 51
rect 355 46 364 48
rect 355 44 360 46
rect 362 44 364 46
rect 355 42 364 44
rect 374 47 380 49
rect 374 45 376 47
rect 378 45 380 47
rect 384 47 386 49
rect 388 47 390 49
rect 414 48 416 52
rect 425 48 427 52
rect 384 45 390 47
rect 374 43 380 45
rect 343 39 345 42
rect 357 39 359 42
rect 375 39 377 43
rect 275 21 277 26
rect 312 21 314 26
rect 133 7 190 9
rect 223 12 225 17
rect 233 9 235 17
rect 243 13 245 17
rect 257 13 259 17
rect 288 9 290 21
rect 388 31 390 45
rect 410 46 416 48
rect 410 44 412 46
rect 414 44 416 46
rect 410 42 416 44
rect 421 46 427 48
rect 435 49 437 52
rect 435 47 449 49
rect 421 44 423 46
rect 425 44 427 46
rect 421 42 427 44
rect 443 46 449 47
rect 443 44 445 46
rect 447 44 449 46
rect 412 39 414 42
rect 423 39 425 42
rect 433 39 435 43
rect 443 42 449 44
rect 455 48 457 54
rect 475 49 477 54
rect 488 51 490 54
rect 555 65 557 69
rect 545 53 547 57
rect 575 64 577 69
rect 588 61 590 73
rect 645 73 690 75
rect 645 68 647 73
rect 614 62 616 66
rect 625 63 627 68
rect 635 63 637 68
rect 484 49 490 51
rect 455 46 464 48
rect 455 44 460 46
rect 462 44 464 46
rect 455 42 464 44
rect 474 47 480 49
rect 474 45 476 47
rect 478 45 480 47
rect 484 47 486 49
rect 488 47 490 49
rect 514 48 516 52
rect 525 48 527 52
rect 484 45 490 47
rect 474 43 480 45
rect 443 39 445 42
rect 457 39 459 42
rect 475 39 477 43
rect 375 21 377 26
rect 412 21 414 26
rect 233 7 290 9
rect 323 12 325 17
rect 333 9 335 17
rect 343 13 345 17
rect 357 13 359 17
rect 388 9 390 21
rect 488 31 490 45
rect 510 46 516 48
rect 510 44 512 46
rect 514 44 516 46
rect 510 42 516 44
rect 521 46 527 48
rect 535 49 537 52
rect 535 47 549 49
rect 521 44 523 46
rect 525 44 527 46
rect 521 42 527 44
rect 543 46 549 47
rect 543 44 545 46
rect 547 44 549 46
rect 512 39 514 42
rect 523 39 525 42
rect 533 39 535 43
rect 543 42 549 44
rect 555 48 557 54
rect 575 49 577 54
rect 588 51 590 54
rect 655 65 657 69
rect 645 53 647 57
rect 675 64 677 69
rect 688 61 690 73
rect 745 73 790 75
rect 745 68 747 73
rect 714 62 716 66
rect 725 63 727 68
rect 735 63 737 68
rect 584 49 590 51
rect 555 46 564 48
rect 555 44 560 46
rect 562 44 564 46
rect 555 42 564 44
rect 574 47 580 49
rect 574 45 576 47
rect 578 45 580 47
rect 584 47 586 49
rect 588 47 590 49
rect 614 48 616 52
rect 625 48 627 52
rect 584 45 590 47
rect 574 43 580 45
rect 543 39 545 42
rect 557 39 559 42
rect 575 39 577 43
rect 475 21 477 26
rect 512 21 514 26
rect 333 7 390 9
rect 423 12 425 17
rect 433 9 435 17
rect 443 13 445 17
rect 457 13 459 17
rect 488 9 490 21
rect 588 31 590 45
rect 610 46 616 48
rect 610 44 612 46
rect 614 44 616 46
rect 610 42 616 44
rect 621 46 627 48
rect 635 49 637 52
rect 635 47 649 49
rect 621 44 623 46
rect 625 44 627 46
rect 621 42 627 44
rect 643 46 649 47
rect 643 44 645 46
rect 647 44 649 46
rect 612 39 614 42
rect 623 39 625 42
rect 633 39 635 43
rect 643 42 649 44
rect 655 48 657 54
rect 675 49 677 54
rect 688 51 690 54
rect 755 65 757 69
rect 745 53 747 57
rect 775 64 777 69
rect 788 61 790 73
rect 684 49 690 51
rect 655 46 664 48
rect 655 44 660 46
rect 662 44 664 46
rect 655 42 664 44
rect 674 47 680 49
rect 674 45 676 47
rect 678 45 680 47
rect 684 47 686 49
rect 688 47 690 49
rect 714 48 716 52
rect 725 48 727 52
rect 684 45 690 47
rect 674 43 680 45
rect 643 39 645 42
rect 657 39 659 42
rect 675 39 677 43
rect 575 21 577 26
rect 612 21 614 26
rect 433 7 490 9
rect 523 12 525 17
rect 533 9 535 17
rect 543 13 545 17
rect 557 13 559 17
rect 588 9 590 21
rect 688 31 690 45
rect 710 46 716 48
rect 710 44 712 46
rect 714 44 716 46
rect 710 42 716 44
rect 721 46 727 48
rect 735 49 737 52
rect 735 47 749 49
rect 721 44 723 46
rect 725 44 727 46
rect 721 42 727 44
rect 743 46 749 47
rect 743 44 745 46
rect 747 44 749 46
rect 712 39 714 42
rect 723 39 725 42
rect 733 39 735 43
rect 743 42 749 44
rect 755 48 757 54
rect 775 49 777 54
rect 788 51 790 54
rect 784 49 790 51
rect 755 46 764 48
rect 755 44 760 46
rect 762 44 764 46
rect 755 42 764 44
rect 774 47 780 49
rect 774 45 776 47
rect 778 45 780 47
rect 784 47 786 49
rect 788 47 790 49
rect 784 45 790 47
rect 774 43 780 45
rect 743 39 745 42
rect 757 39 759 42
rect 775 39 777 43
rect 675 21 677 26
rect 712 21 714 26
rect 533 7 590 9
rect 623 12 625 17
rect 633 9 635 17
rect 643 13 645 17
rect 657 13 659 17
rect 688 9 690 21
rect 788 31 790 45
rect 775 21 777 26
rect 633 7 690 9
rect 723 12 725 17
rect 733 9 735 17
rect 743 13 745 17
rect 757 13 759 17
rect 788 9 790 21
rect 733 7 790 9
rect 16 -27 73 -25
rect 6 -35 8 -30
rect 16 -35 18 -27
rect 26 -35 28 -31
rect 40 -35 42 -31
rect -5 -44 -3 -39
rect 71 -39 73 -27
rect 122 -27 179 -25
rect 112 -35 114 -30
rect 122 -35 124 -27
rect 132 -35 134 -31
rect 146 -35 148 -31
rect 58 -44 60 -39
rect 101 -44 103 -39
rect -5 -60 -3 -57
rect 6 -60 8 -57
rect -7 -62 -1 -60
rect -7 -64 -5 -62
rect -3 -64 -1 -62
rect -7 -66 -1 -64
rect 4 -62 10 -60
rect 16 -61 18 -57
rect 26 -60 28 -57
rect 40 -60 42 -57
rect 4 -64 6 -62
rect 8 -64 10 -62
rect 4 -66 10 -64
rect 26 -62 32 -60
rect 26 -64 28 -62
rect 30 -64 32 -62
rect 26 -65 32 -64
rect -3 -70 -1 -66
rect 8 -70 10 -66
rect 18 -67 32 -65
rect 38 -62 47 -60
rect 58 -61 60 -57
rect 38 -64 43 -62
rect 45 -64 47 -62
rect 38 -66 47 -64
rect 57 -63 63 -61
rect 71 -63 73 -49
rect 177 -39 179 -27
rect 228 -27 285 -25
rect 218 -35 220 -30
rect 228 -35 230 -27
rect 238 -35 240 -31
rect 252 -35 254 -31
rect 164 -44 166 -39
rect 207 -44 209 -39
rect 101 -60 103 -57
rect 112 -60 114 -57
rect 57 -65 59 -63
rect 61 -65 63 -63
rect 18 -70 20 -67
rect -3 -84 -1 -80
rect 28 -75 30 -71
rect 38 -72 40 -66
rect 57 -67 63 -65
rect 67 -65 73 -63
rect 67 -67 69 -65
rect 71 -67 73 -65
rect 99 -62 105 -60
rect 99 -64 101 -62
rect 103 -64 105 -62
rect 99 -66 105 -64
rect 110 -62 116 -60
rect 122 -61 124 -57
rect 132 -60 134 -57
rect 146 -60 148 -57
rect 110 -64 112 -62
rect 114 -64 116 -62
rect 110 -66 116 -64
rect 132 -62 138 -60
rect 132 -64 134 -62
rect 136 -64 138 -62
rect 132 -65 138 -64
rect 58 -72 60 -67
rect 67 -69 73 -67
rect 71 -72 73 -69
rect 103 -70 105 -66
rect 114 -70 116 -66
rect 124 -67 138 -65
rect 144 -62 153 -60
rect 164 -61 166 -57
rect 144 -64 149 -62
rect 151 -64 153 -62
rect 144 -66 153 -64
rect 163 -63 169 -61
rect 177 -63 179 -49
rect 283 -39 285 -27
rect 334 -27 391 -25
rect 324 -35 326 -30
rect 334 -35 336 -27
rect 344 -35 346 -31
rect 358 -35 360 -31
rect 270 -44 272 -39
rect 313 -44 315 -39
rect 207 -60 209 -57
rect 218 -60 220 -57
rect 163 -65 165 -63
rect 167 -65 169 -63
rect 124 -70 126 -67
rect 8 -86 10 -81
rect 18 -86 20 -81
rect 28 -91 30 -86
rect 38 -87 40 -83
rect 58 -87 60 -82
rect 71 -91 73 -79
rect 103 -84 105 -80
rect 134 -75 136 -71
rect 144 -72 146 -66
rect 163 -67 169 -65
rect 173 -65 179 -63
rect 173 -67 175 -65
rect 177 -67 179 -65
rect 205 -62 211 -60
rect 205 -64 207 -62
rect 209 -64 211 -62
rect 205 -66 211 -64
rect 216 -62 222 -60
rect 228 -61 230 -57
rect 238 -60 240 -57
rect 252 -60 254 -57
rect 216 -64 218 -62
rect 220 -64 222 -62
rect 216 -66 222 -64
rect 238 -62 244 -60
rect 238 -64 240 -62
rect 242 -64 244 -62
rect 238 -65 244 -64
rect 164 -72 166 -67
rect 173 -69 179 -67
rect 177 -72 179 -69
rect 209 -70 211 -66
rect 220 -70 222 -66
rect 230 -67 244 -65
rect 250 -62 259 -60
rect 270 -61 272 -57
rect 250 -64 255 -62
rect 257 -64 259 -62
rect 250 -66 259 -64
rect 269 -63 275 -61
rect 283 -63 285 -49
rect 389 -39 391 -27
rect 440 -27 497 -25
rect 430 -35 432 -30
rect 440 -35 442 -27
rect 450 -35 452 -31
rect 464 -35 466 -31
rect 376 -44 378 -39
rect 419 -44 421 -39
rect 313 -60 315 -57
rect 324 -60 326 -57
rect 269 -65 271 -63
rect 273 -65 275 -63
rect 230 -70 232 -67
rect 114 -86 116 -81
rect 124 -86 126 -81
rect 28 -93 73 -91
rect 134 -91 136 -86
rect 144 -87 146 -83
rect 164 -87 166 -82
rect 177 -91 179 -79
rect 209 -84 211 -80
rect 240 -75 242 -71
rect 250 -72 252 -66
rect 269 -67 275 -65
rect 279 -65 285 -63
rect 279 -67 281 -65
rect 283 -67 285 -65
rect 311 -62 317 -60
rect 311 -64 313 -62
rect 315 -64 317 -62
rect 311 -66 317 -64
rect 322 -62 328 -60
rect 334 -61 336 -57
rect 344 -60 346 -57
rect 358 -60 360 -57
rect 322 -64 324 -62
rect 326 -64 328 -62
rect 322 -66 328 -64
rect 344 -62 350 -60
rect 344 -64 346 -62
rect 348 -64 350 -62
rect 344 -65 350 -64
rect 270 -72 272 -67
rect 279 -69 285 -67
rect 283 -72 285 -69
rect 315 -70 317 -66
rect 326 -70 328 -66
rect 336 -67 350 -65
rect 356 -62 365 -60
rect 376 -61 378 -57
rect 356 -64 361 -62
rect 363 -64 365 -62
rect 356 -66 365 -64
rect 375 -63 381 -61
rect 389 -63 391 -49
rect 495 -39 497 -27
rect 546 -27 603 -25
rect 536 -35 538 -30
rect 546 -35 548 -27
rect 556 -35 558 -31
rect 570 -35 572 -31
rect 482 -44 484 -39
rect 525 -44 527 -39
rect 419 -60 421 -57
rect 430 -60 432 -57
rect 375 -65 377 -63
rect 379 -65 381 -63
rect 336 -70 338 -67
rect 220 -86 222 -81
rect 230 -86 232 -81
rect 134 -93 179 -91
rect 240 -91 242 -86
rect 250 -87 252 -83
rect 270 -87 272 -82
rect 283 -91 285 -79
rect 315 -84 317 -80
rect 346 -75 348 -71
rect 356 -72 358 -66
rect 375 -67 381 -65
rect 385 -65 391 -63
rect 385 -67 387 -65
rect 389 -67 391 -65
rect 417 -62 423 -60
rect 417 -64 419 -62
rect 421 -64 423 -62
rect 417 -66 423 -64
rect 428 -62 434 -60
rect 440 -61 442 -57
rect 450 -60 452 -57
rect 464 -60 466 -57
rect 428 -64 430 -62
rect 432 -64 434 -62
rect 428 -66 434 -64
rect 450 -62 456 -60
rect 450 -64 452 -62
rect 454 -64 456 -62
rect 450 -65 456 -64
rect 376 -72 378 -67
rect 385 -69 391 -67
rect 389 -72 391 -69
rect 421 -70 423 -66
rect 432 -70 434 -66
rect 442 -67 456 -65
rect 462 -62 471 -60
rect 482 -61 484 -57
rect 462 -64 467 -62
rect 469 -64 471 -62
rect 462 -66 471 -64
rect 481 -63 487 -61
rect 495 -63 497 -49
rect 601 -39 603 -27
rect 652 -27 709 -25
rect 642 -35 644 -30
rect 652 -35 654 -27
rect 662 -35 664 -31
rect 676 -35 678 -31
rect 588 -44 590 -39
rect 631 -44 633 -39
rect 525 -60 527 -57
rect 536 -60 538 -57
rect 481 -65 483 -63
rect 485 -65 487 -63
rect 442 -70 444 -67
rect 326 -86 328 -81
rect 336 -86 338 -81
rect 240 -93 285 -91
rect 346 -91 348 -86
rect 356 -87 358 -83
rect 376 -87 378 -82
rect 389 -91 391 -79
rect 421 -84 423 -80
rect 452 -75 454 -71
rect 462 -72 464 -66
rect 481 -67 487 -65
rect 491 -65 497 -63
rect 491 -67 493 -65
rect 495 -67 497 -65
rect 523 -62 529 -60
rect 523 -64 525 -62
rect 527 -64 529 -62
rect 523 -66 529 -64
rect 534 -62 540 -60
rect 546 -61 548 -57
rect 556 -60 558 -57
rect 570 -60 572 -57
rect 534 -64 536 -62
rect 538 -64 540 -62
rect 534 -66 540 -64
rect 556 -62 562 -60
rect 556 -64 558 -62
rect 560 -64 562 -62
rect 556 -65 562 -64
rect 482 -72 484 -67
rect 491 -69 497 -67
rect 495 -72 497 -69
rect 527 -70 529 -66
rect 538 -70 540 -66
rect 548 -67 562 -65
rect 568 -62 577 -60
rect 588 -61 590 -57
rect 568 -64 573 -62
rect 575 -64 577 -62
rect 568 -66 577 -64
rect 587 -63 593 -61
rect 601 -63 603 -49
rect 707 -39 709 -27
rect 758 -27 815 -25
rect 748 -35 750 -30
rect 758 -35 760 -27
rect 768 -35 770 -31
rect 782 -35 784 -31
rect 694 -44 696 -39
rect 737 -44 739 -39
rect 631 -60 633 -57
rect 642 -60 644 -57
rect 587 -65 589 -63
rect 591 -65 593 -63
rect 548 -70 550 -67
rect 432 -86 434 -81
rect 442 -86 444 -81
rect 346 -93 391 -91
rect 452 -91 454 -86
rect 462 -87 464 -83
rect 482 -87 484 -82
rect 495 -91 497 -79
rect 527 -84 529 -80
rect 558 -75 560 -71
rect 568 -72 570 -66
rect 587 -67 593 -65
rect 597 -65 603 -63
rect 597 -67 599 -65
rect 601 -67 603 -65
rect 629 -62 635 -60
rect 629 -64 631 -62
rect 633 -64 635 -62
rect 629 -66 635 -64
rect 640 -62 646 -60
rect 652 -61 654 -57
rect 662 -60 664 -57
rect 676 -60 678 -57
rect 640 -64 642 -62
rect 644 -64 646 -62
rect 640 -66 646 -64
rect 662 -62 668 -60
rect 662 -64 664 -62
rect 666 -64 668 -62
rect 662 -65 668 -64
rect 588 -72 590 -67
rect 597 -69 603 -67
rect 601 -72 603 -69
rect 633 -70 635 -66
rect 644 -70 646 -66
rect 654 -67 668 -65
rect 674 -62 683 -60
rect 694 -61 696 -57
rect 674 -64 679 -62
rect 681 -64 683 -62
rect 674 -66 683 -64
rect 693 -63 699 -61
rect 707 -63 709 -49
rect 813 -39 815 -27
rect 864 -27 921 -25
rect 854 -35 856 -30
rect 864 -35 866 -27
rect 874 -35 876 -31
rect 888 -35 890 -31
rect 800 -44 802 -39
rect 843 -44 845 -39
rect 737 -60 739 -57
rect 748 -60 750 -57
rect 693 -65 695 -63
rect 697 -65 699 -63
rect 654 -70 656 -67
rect 538 -86 540 -81
rect 548 -86 550 -81
rect 452 -93 497 -91
rect 558 -91 560 -86
rect 568 -87 570 -83
rect 588 -87 590 -82
rect 601 -91 603 -79
rect 633 -84 635 -80
rect 664 -75 666 -71
rect 674 -72 676 -66
rect 693 -67 699 -65
rect 703 -65 709 -63
rect 703 -67 705 -65
rect 707 -67 709 -65
rect 735 -62 741 -60
rect 735 -64 737 -62
rect 739 -64 741 -62
rect 735 -66 741 -64
rect 746 -62 752 -60
rect 758 -61 760 -57
rect 768 -60 770 -57
rect 782 -60 784 -57
rect 746 -64 748 -62
rect 750 -64 752 -62
rect 746 -66 752 -64
rect 768 -62 774 -60
rect 768 -64 770 -62
rect 772 -64 774 -62
rect 768 -65 774 -64
rect 694 -72 696 -67
rect 703 -69 709 -67
rect 707 -72 709 -69
rect 739 -70 741 -66
rect 750 -70 752 -66
rect 760 -67 774 -65
rect 780 -62 789 -60
rect 800 -61 802 -57
rect 780 -64 785 -62
rect 787 -64 789 -62
rect 780 -66 789 -64
rect 799 -63 805 -61
rect 813 -63 815 -49
rect 919 -39 921 -27
rect 906 -44 908 -39
rect 843 -60 845 -57
rect 854 -60 856 -57
rect 799 -65 801 -63
rect 803 -65 805 -63
rect 760 -70 762 -67
rect 644 -86 646 -81
rect 654 -86 656 -81
rect 558 -93 603 -91
rect 664 -91 666 -86
rect 674 -87 676 -83
rect 694 -87 696 -82
rect 707 -91 709 -79
rect 739 -84 741 -80
rect 770 -75 772 -71
rect 780 -72 782 -66
rect 799 -67 805 -65
rect 809 -65 815 -63
rect 809 -67 811 -65
rect 813 -67 815 -65
rect 841 -62 847 -60
rect 841 -64 843 -62
rect 845 -64 847 -62
rect 841 -66 847 -64
rect 852 -62 858 -60
rect 864 -61 866 -57
rect 874 -60 876 -57
rect 888 -60 890 -57
rect 852 -64 854 -62
rect 856 -64 858 -62
rect 852 -66 858 -64
rect 874 -62 880 -60
rect 874 -64 876 -62
rect 878 -64 880 -62
rect 874 -65 880 -64
rect 800 -72 802 -67
rect 809 -69 815 -67
rect 813 -72 815 -69
rect 845 -70 847 -66
rect 856 -70 858 -66
rect 866 -67 880 -65
rect 886 -62 895 -60
rect 906 -61 908 -57
rect 886 -64 891 -62
rect 893 -64 895 -62
rect 886 -66 895 -64
rect 905 -63 911 -61
rect 919 -63 921 -49
rect 905 -65 907 -63
rect 909 -65 911 -63
rect 866 -70 868 -67
rect 750 -86 752 -81
rect 760 -86 762 -81
rect 664 -93 709 -91
rect 770 -91 772 -86
rect 780 -87 782 -83
rect 800 -87 802 -82
rect 813 -91 815 -79
rect 845 -84 847 -80
rect 876 -75 878 -71
rect 886 -72 888 -66
rect 905 -67 911 -65
rect 915 -65 921 -63
rect 915 -67 917 -65
rect 919 -67 921 -65
rect 906 -72 908 -67
rect 915 -69 921 -67
rect 919 -72 921 -69
rect 856 -86 858 -81
rect 866 -86 868 -81
rect 770 -93 815 -91
rect 876 -91 878 -86
rect 886 -87 888 -83
rect 906 -87 908 -82
rect 919 -91 921 -79
rect 876 -93 921 -91
<< ndif >>
rect 134 1183 140 1185
rect 134 1181 136 1183
rect 138 1181 140 1183
rect 134 1179 140 1181
rect 118 1176 123 1179
rect 94 1174 103 1176
rect 94 1172 96 1174
rect 98 1172 103 1174
rect 94 1171 103 1172
rect 82 1168 87 1171
rect 80 1166 87 1168
rect 80 1164 82 1166
rect 84 1164 87 1166
rect 80 1162 87 1164
rect 89 1167 103 1171
rect 105 1171 113 1176
rect 105 1169 108 1171
rect 110 1169 113 1171
rect 105 1167 113 1169
rect 115 1173 123 1176
rect 115 1171 118 1173
rect 120 1171 123 1173
rect 115 1167 123 1171
rect 125 1167 130 1179
rect 132 1167 140 1179
rect 148 1183 154 1185
rect 148 1181 150 1183
rect 152 1181 154 1183
rect 148 1176 154 1181
rect 195 1183 202 1185
rect 195 1181 197 1183
rect 199 1181 202 1183
rect 148 1168 156 1176
rect 158 1174 165 1176
rect 158 1172 161 1174
rect 163 1173 165 1174
rect 195 1175 202 1181
rect 282 1183 288 1185
rect 282 1181 284 1183
rect 286 1181 288 1183
rect 336 1183 343 1185
rect 336 1182 338 1183
rect 282 1179 288 1181
rect 266 1176 271 1179
rect 195 1173 204 1175
rect 163 1172 167 1173
rect 158 1168 167 1172
rect 89 1162 94 1167
rect 162 1165 167 1168
rect 169 1171 176 1173
rect 169 1169 172 1171
rect 174 1169 176 1171
rect 169 1165 176 1169
rect 184 1171 191 1173
rect 184 1169 186 1171
rect 188 1169 191 1171
rect 184 1167 191 1169
rect 186 1164 191 1167
rect 193 1164 204 1173
rect 206 1164 211 1175
rect 213 1173 220 1175
rect 213 1171 216 1173
rect 218 1171 220 1173
rect 242 1174 251 1176
rect 242 1172 244 1174
rect 246 1172 251 1174
rect 242 1171 251 1172
rect 213 1169 220 1171
rect 213 1164 218 1169
rect 230 1168 235 1171
rect 228 1166 235 1168
rect 228 1164 230 1166
rect 232 1164 235 1166
rect 228 1162 235 1164
rect 237 1167 251 1171
rect 253 1171 261 1176
rect 253 1169 256 1171
rect 258 1169 261 1171
rect 253 1167 261 1169
rect 263 1173 271 1176
rect 263 1171 266 1173
rect 268 1171 271 1173
rect 263 1167 271 1171
rect 273 1167 278 1179
rect 280 1167 288 1179
rect 306 1176 311 1182
rect 304 1174 311 1176
rect 304 1172 306 1174
rect 308 1172 311 1174
rect 304 1170 311 1172
rect 237 1162 242 1167
rect 306 1162 311 1170
rect 313 1162 318 1182
rect 320 1162 325 1182
rect 327 1162 332 1182
rect 334 1181 338 1182
rect 340 1181 343 1183
rect 334 1162 343 1181
rect 566 1173 572 1175
rect 566 1171 568 1173
rect 570 1172 572 1173
rect 658 1183 664 1185
rect 658 1181 660 1183
rect 662 1181 664 1183
rect 658 1179 664 1181
rect 642 1176 647 1179
rect 618 1174 627 1176
rect 570 1171 574 1172
rect 360 1168 365 1171
rect 358 1166 365 1168
rect 358 1164 360 1166
rect 362 1164 365 1166
rect 358 1162 365 1164
rect 367 1169 378 1171
rect 367 1167 374 1169
rect 376 1167 378 1169
rect 367 1162 378 1167
rect 566 1162 574 1171
rect 576 1166 584 1172
rect 576 1164 579 1166
rect 581 1164 584 1166
rect 576 1162 584 1164
rect 586 1170 594 1172
rect 618 1172 620 1174
rect 622 1172 627 1174
rect 618 1171 627 1172
rect 586 1168 590 1170
rect 592 1168 594 1170
rect 606 1168 611 1171
rect 586 1162 594 1168
rect 604 1166 611 1168
rect 604 1164 606 1166
rect 608 1164 611 1166
rect 604 1162 611 1164
rect 613 1167 627 1171
rect 629 1171 637 1176
rect 629 1169 632 1171
rect 634 1169 637 1171
rect 629 1167 637 1169
rect 639 1173 647 1176
rect 639 1171 642 1173
rect 644 1171 647 1173
rect 639 1167 647 1171
rect 649 1167 654 1179
rect 656 1167 664 1179
rect 677 1168 682 1171
rect 613 1162 618 1167
rect 675 1166 682 1168
rect 675 1164 677 1166
rect 679 1164 682 1166
rect 675 1162 682 1164
rect 684 1169 695 1171
rect 714 1180 722 1182
rect 714 1178 717 1180
rect 719 1178 722 1180
rect 714 1173 722 1178
rect 714 1171 717 1173
rect 719 1171 722 1173
rect 684 1167 691 1169
rect 693 1167 695 1169
rect 714 1167 722 1171
rect 724 1173 732 1182
rect 724 1171 727 1173
rect 729 1171 732 1173
rect 724 1167 732 1171
rect 734 1180 742 1182
rect 734 1178 737 1180
rect 739 1178 742 1180
rect 734 1167 742 1178
rect 684 1162 695 1167
rect 85 1062 90 1070
rect 83 1060 90 1062
rect 83 1058 85 1060
rect 87 1058 90 1060
rect 83 1056 90 1058
rect 85 1050 90 1056
rect 92 1050 97 1070
rect 99 1061 108 1070
rect 116 1068 123 1070
rect 116 1066 118 1068
rect 120 1066 123 1068
rect 116 1064 123 1066
rect 118 1061 123 1064
rect 125 1065 136 1070
rect 146 1065 151 1068
rect 125 1063 132 1065
rect 134 1063 136 1065
rect 125 1061 136 1063
rect 144 1063 151 1065
rect 144 1061 146 1063
rect 148 1061 151 1063
rect 99 1059 104 1061
rect 106 1059 108 1061
rect 99 1054 108 1059
rect 144 1059 151 1061
rect 153 1059 164 1068
rect 155 1057 164 1059
rect 166 1057 171 1068
rect 173 1063 178 1068
rect 188 1067 195 1069
rect 188 1065 190 1067
rect 192 1065 195 1067
rect 188 1063 195 1065
rect 173 1061 180 1063
rect 173 1059 176 1061
rect 178 1059 180 1061
rect 190 1060 195 1063
rect 197 1060 208 1069
rect 173 1057 180 1059
rect 99 1052 104 1054
rect 106 1052 108 1054
rect 99 1050 108 1052
rect 155 1051 162 1057
rect 199 1056 208 1060
rect 210 1056 215 1069
rect 217 1056 222 1069
rect 224 1062 229 1069
rect 224 1060 231 1062
rect 224 1058 227 1060
rect 229 1058 231 1060
rect 224 1056 231 1058
rect 256 1060 263 1062
rect 256 1058 258 1060
rect 260 1058 263 1060
rect 256 1056 263 1058
rect 265 1060 273 1062
rect 265 1058 268 1060
rect 270 1058 273 1060
rect 265 1056 273 1058
rect 275 1056 285 1062
rect 287 1060 295 1062
rect 287 1058 290 1060
rect 292 1058 295 1060
rect 287 1056 295 1058
rect 297 1060 304 1062
rect 297 1058 300 1060
rect 302 1058 304 1060
rect 297 1056 304 1058
rect 155 1049 157 1051
rect 159 1049 162 1051
rect 155 1047 162 1049
rect 199 1051 206 1056
rect 277 1051 283 1056
rect 569 1065 580 1070
rect 569 1063 571 1065
rect 573 1063 580 1065
rect 569 1061 580 1063
rect 582 1068 589 1070
rect 582 1066 585 1068
rect 587 1066 589 1068
rect 582 1064 589 1066
rect 603 1065 608 1068
rect 582 1061 587 1064
rect 601 1063 608 1065
rect 601 1061 603 1063
rect 605 1061 608 1063
rect 601 1059 608 1061
rect 610 1059 621 1068
rect 612 1057 621 1059
rect 623 1057 628 1068
rect 630 1063 635 1068
rect 630 1061 637 1063
rect 630 1059 633 1061
rect 635 1059 637 1061
rect 630 1057 637 1059
rect 647 1061 656 1070
rect 647 1059 649 1061
rect 651 1059 656 1061
rect 199 1049 201 1051
rect 203 1049 206 1051
rect 199 1047 206 1049
rect 277 1049 279 1051
rect 281 1049 283 1051
rect 277 1047 283 1049
rect 612 1051 619 1057
rect 647 1054 656 1059
rect 647 1052 649 1054
rect 651 1052 656 1054
rect 612 1049 614 1051
rect 616 1049 619 1051
rect 647 1050 656 1052
rect 658 1050 663 1070
rect 665 1062 670 1070
rect 729 1065 734 1070
rect 665 1060 672 1062
rect 665 1058 668 1060
rect 670 1058 672 1060
rect 665 1056 672 1058
rect 665 1050 670 1056
rect 683 1053 691 1065
rect 693 1053 698 1065
rect 700 1061 708 1065
rect 700 1059 703 1061
rect 705 1059 708 1061
rect 700 1056 708 1059
rect 710 1063 718 1065
rect 710 1061 713 1063
rect 715 1061 718 1063
rect 710 1056 718 1061
rect 720 1061 734 1065
rect 736 1068 743 1070
rect 736 1066 739 1068
rect 741 1066 743 1068
rect 736 1064 743 1066
rect 736 1061 741 1064
rect 720 1060 729 1061
rect 720 1058 725 1060
rect 727 1058 729 1060
rect 720 1056 729 1058
rect 700 1053 705 1056
rect 683 1051 689 1053
rect 612 1047 619 1049
rect 683 1049 685 1051
rect 687 1049 689 1051
rect 683 1047 689 1049
rect 134 1039 140 1041
rect 134 1037 136 1039
rect 138 1037 140 1039
rect 134 1035 140 1037
rect 118 1032 123 1035
rect 94 1030 103 1032
rect 94 1028 96 1030
rect 98 1028 103 1030
rect 94 1027 103 1028
rect 82 1024 87 1027
rect 80 1022 87 1024
rect 80 1020 82 1022
rect 84 1020 87 1022
rect 80 1018 87 1020
rect 89 1023 103 1027
rect 105 1027 113 1032
rect 105 1025 108 1027
rect 110 1025 113 1027
rect 105 1023 113 1025
rect 115 1029 123 1032
rect 115 1027 118 1029
rect 120 1027 123 1029
rect 115 1023 123 1027
rect 125 1023 130 1035
rect 132 1023 140 1035
rect 153 1032 158 1038
rect 151 1030 158 1032
rect 151 1028 153 1030
rect 155 1028 158 1030
rect 151 1026 158 1028
rect 89 1018 94 1023
rect 153 1018 158 1026
rect 160 1018 165 1038
rect 167 1036 176 1038
rect 167 1034 172 1036
rect 174 1034 176 1036
rect 167 1029 176 1034
rect 167 1027 172 1029
rect 174 1027 176 1029
rect 167 1018 176 1027
rect 208 1039 215 1041
rect 208 1037 211 1039
rect 213 1037 215 1039
rect 208 1036 215 1037
rect 231 1039 237 1041
rect 231 1037 233 1039
rect 235 1037 237 1039
rect 231 1036 237 1037
rect 290 1039 297 1041
rect 290 1037 293 1039
rect 295 1037 297 1039
rect 208 1026 217 1036
rect 219 1030 227 1036
rect 219 1028 222 1030
rect 224 1028 227 1030
rect 219 1026 227 1028
rect 229 1026 239 1036
rect 241 1032 246 1036
rect 290 1032 297 1037
rect 645 1039 652 1041
rect 241 1030 248 1032
rect 241 1028 244 1030
rect 246 1028 248 1030
rect 241 1026 248 1028
rect 265 1030 272 1032
rect 265 1028 267 1030
rect 269 1028 272 1030
rect 265 1026 272 1028
rect 267 1019 272 1026
rect 274 1019 279 1032
rect 281 1019 286 1032
rect 288 1028 297 1032
rect 288 1019 299 1028
rect 301 1025 306 1028
rect 301 1023 308 1025
rect 513 1024 518 1027
rect 301 1021 304 1023
rect 306 1021 308 1023
rect 301 1019 308 1021
rect 511 1022 518 1024
rect 511 1020 513 1022
rect 515 1020 518 1022
rect 511 1018 518 1020
rect 520 1025 531 1027
rect 590 1036 598 1038
rect 590 1034 593 1036
rect 595 1034 598 1036
rect 590 1029 598 1034
rect 590 1027 593 1029
rect 595 1027 598 1029
rect 520 1023 527 1025
rect 529 1023 531 1025
rect 590 1023 598 1027
rect 600 1029 608 1038
rect 600 1027 603 1029
rect 605 1027 608 1029
rect 600 1023 608 1027
rect 610 1036 618 1038
rect 645 1037 648 1039
rect 650 1037 652 1039
rect 610 1034 613 1036
rect 615 1034 618 1036
rect 610 1023 618 1034
rect 645 1031 652 1037
rect 627 1029 634 1031
rect 627 1027 629 1029
rect 631 1027 634 1029
rect 627 1025 634 1027
rect 520 1018 531 1023
rect 629 1020 634 1025
rect 636 1020 641 1031
rect 643 1029 652 1031
rect 643 1020 654 1029
rect 656 1027 663 1029
rect 656 1025 659 1027
rect 661 1025 663 1027
rect 656 1023 663 1025
rect 675 1024 680 1027
rect 656 1020 661 1023
rect 673 1022 680 1024
rect 673 1020 675 1022
rect 677 1020 680 1022
rect 673 1018 680 1020
rect 682 1025 693 1027
rect 714 1036 722 1038
rect 714 1034 717 1036
rect 719 1034 722 1036
rect 714 1029 722 1034
rect 714 1027 717 1029
rect 719 1027 722 1029
rect 682 1023 689 1025
rect 691 1023 693 1025
rect 714 1023 722 1027
rect 724 1029 732 1038
rect 724 1027 727 1029
rect 729 1027 732 1029
rect 724 1023 732 1027
rect 734 1036 742 1038
rect 734 1034 737 1036
rect 739 1034 742 1036
rect 734 1023 742 1034
rect 682 1018 693 1023
rect 116 924 123 926
rect 94 920 99 923
rect 80 917 88 920
rect 77 913 88 917
rect 80 912 88 913
rect 90 916 99 920
rect 90 914 93 916
rect 95 915 99 916
rect 101 919 108 923
rect 116 922 118 924
rect 120 922 123 924
rect 116 920 123 922
rect 101 917 104 919
rect 106 917 108 919
rect 118 917 123 920
rect 125 921 136 926
rect 146 921 151 924
rect 125 919 132 921
rect 134 919 136 921
rect 125 917 136 919
rect 144 919 151 921
rect 144 917 146 919
rect 148 917 151 919
rect 101 915 108 917
rect 95 914 97 915
rect 90 912 97 914
rect 80 907 86 912
rect 144 915 151 917
rect 153 915 164 924
rect 155 913 164 915
rect 166 913 171 924
rect 173 919 178 924
rect 246 921 251 926
rect 173 917 180 919
rect 173 915 176 917
rect 178 915 180 917
rect 173 913 180 915
rect 80 905 82 907
rect 84 905 86 907
rect 80 903 86 905
rect 155 907 162 913
rect 200 909 208 921
rect 210 909 215 921
rect 217 917 225 921
rect 217 915 220 917
rect 222 915 225 917
rect 217 912 225 915
rect 227 919 235 921
rect 227 917 230 919
rect 232 917 235 919
rect 227 912 235 917
rect 237 917 251 921
rect 253 924 260 926
rect 253 922 256 924
rect 258 922 260 924
rect 253 920 260 922
rect 253 917 258 920
rect 270 919 275 924
rect 268 917 275 919
rect 237 916 246 917
rect 237 914 242 916
rect 244 914 246 916
rect 237 912 246 914
rect 268 915 270 917
rect 272 915 275 917
rect 268 913 275 915
rect 277 913 282 924
rect 284 915 295 924
rect 297 921 302 924
rect 557 921 562 926
rect 297 919 304 921
rect 297 917 300 919
rect 302 917 304 919
rect 297 915 304 917
rect 284 913 293 915
rect 217 909 222 912
rect 155 905 157 907
rect 159 905 162 907
rect 155 903 162 905
rect 200 907 206 909
rect 200 905 202 907
rect 204 905 206 907
rect 200 903 206 905
rect 286 907 293 913
rect 511 909 519 921
rect 521 909 526 921
rect 528 917 536 921
rect 528 915 531 917
rect 533 915 536 917
rect 528 912 536 915
rect 538 919 546 921
rect 538 917 541 919
rect 543 917 546 919
rect 538 912 546 917
rect 548 917 562 921
rect 564 924 571 926
rect 623 924 630 926
rect 564 922 567 924
rect 569 922 571 924
rect 564 920 571 922
rect 581 921 586 924
rect 564 917 569 920
rect 579 919 586 921
rect 579 917 581 919
rect 583 917 586 919
rect 548 916 557 917
rect 548 914 553 916
rect 555 914 557 916
rect 579 915 586 917
rect 588 915 599 924
rect 548 912 557 914
rect 528 909 533 912
rect 286 905 289 907
rect 291 905 293 907
rect 286 903 293 905
rect 511 907 517 909
rect 511 905 513 907
rect 515 905 517 907
rect 511 903 517 905
rect 590 913 599 915
rect 601 913 606 924
rect 608 919 613 924
rect 623 922 625 924
rect 627 922 630 924
rect 623 920 630 922
rect 608 917 615 919
rect 608 915 611 917
rect 613 915 615 917
rect 625 915 630 920
rect 632 915 641 926
rect 608 913 615 915
rect 590 907 597 913
rect 634 913 636 915
rect 638 913 641 915
rect 590 905 592 907
rect 594 905 597 907
rect 590 903 597 905
rect 634 907 641 913
rect 643 923 651 926
rect 643 921 646 923
rect 648 921 651 923
rect 643 916 651 921
rect 643 914 646 916
rect 648 914 651 916
rect 643 911 651 914
rect 653 924 661 926
rect 653 922 656 924
rect 658 922 661 924
rect 653 911 661 922
rect 663 918 668 926
rect 729 921 734 926
rect 663 916 670 918
rect 663 914 666 916
rect 668 914 670 916
rect 663 911 670 914
rect 643 907 648 911
rect 683 909 691 921
rect 693 909 698 921
rect 700 917 708 921
rect 700 915 703 917
rect 705 915 708 917
rect 700 912 708 915
rect 710 919 718 921
rect 710 917 713 919
rect 715 917 718 919
rect 710 912 718 917
rect 720 917 734 921
rect 736 924 743 926
rect 736 922 739 924
rect 741 922 743 924
rect 736 920 743 922
rect 736 917 741 920
rect 720 916 729 917
rect 720 914 725 916
rect 727 914 729 916
rect 720 912 729 914
rect 700 909 705 912
rect 683 907 689 909
rect 683 905 685 907
rect 687 905 689 907
rect 683 903 689 905
rect 81 891 93 893
rect 81 889 83 891
rect 85 889 93 891
rect 81 881 93 889
rect 95 881 100 893
rect 102 887 107 893
rect 127 895 134 897
rect 127 893 129 895
rect 131 893 134 895
rect 102 885 109 887
rect 127 887 134 893
rect 176 895 183 897
rect 176 893 178 895
rect 180 893 183 895
rect 127 885 136 887
rect 102 883 105 885
rect 107 883 109 885
rect 102 881 109 883
rect 116 883 123 885
rect 116 881 118 883
rect 120 881 123 883
rect 116 879 123 881
rect 118 876 123 879
rect 125 876 136 885
rect 138 876 143 887
rect 145 885 152 887
rect 176 887 183 893
rect 236 895 243 897
rect 236 893 239 895
rect 241 893 243 895
rect 236 887 243 893
rect 303 895 310 897
rect 303 893 305 895
rect 307 893 310 895
rect 176 885 185 887
rect 145 883 148 885
rect 150 883 152 885
rect 145 881 152 883
rect 165 883 172 885
rect 165 881 167 883
rect 169 881 172 883
rect 145 876 150 881
rect 165 879 172 881
rect 167 876 172 879
rect 174 876 185 885
rect 187 876 192 887
rect 194 885 201 887
rect 194 883 197 885
rect 199 883 201 885
rect 194 881 201 883
rect 218 885 225 887
rect 218 883 220 885
rect 222 883 225 885
rect 218 881 225 883
rect 194 876 199 881
rect 220 876 225 881
rect 227 876 232 887
rect 234 885 243 887
rect 234 876 245 885
rect 247 883 254 885
rect 303 887 310 893
rect 347 895 354 897
rect 347 893 349 895
rect 351 893 354 895
rect 504 895 511 897
rect 504 893 507 895
rect 509 893 511 895
rect 303 885 312 887
rect 292 883 299 885
rect 247 881 250 883
rect 252 881 254 883
rect 247 879 254 881
rect 266 880 271 883
rect 247 876 252 879
rect 264 878 271 880
rect 264 876 266 878
rect 268 876 271 878
rect 264 874 271 876
rect 273 881 284 883
rect 273 879 280 881
rect 282 879 284 881
rect 292 881 294 883
rect 296 881 299 883
rect 292 879 299 881
rect 273 874 284 879
rect 294 876 299 879
rect 301 876 312 885
rect 314 876 319 887
rect 321 885 328 887
rect 321 883 324 885
rect 326 883 328 885
rect 347 888 354 893
rect 347 884 356 888
rect 321 881 328 883
rect 338 881 343 884
rect 321 876 326 881
rect 336 879 343 881
rect 336 877 338 879
rect 340 877 343 879
rect 336 875 343 877
rect 345 875 356 884
rect 358 875 363 888
rect 365 875 370 888
rect 372 886 379 888
rect 504 887 511 893
rect 577 895 584 897
rect 577 893 580 895
rect 582 893 584 895
rect 372 884 375 886
rect 377 884 379 886
rect 372 882 379 884
rect 486 885 493 887
rect 486 883 488 885
rect 490 883 493 885
rect 372 875 377 882
rect 486 881 493 883
rect 488 876 493 881
rect 495 876 500 887
rect 502 885 511 887
rect 502 876 513 885
rect 515 883 522 885
rect 577 887 584 893
rect 618 895 625 897
rect 618 893 620 895
rect 622 893 625 895
rect 681 895 688 897
rect 681 893 684 895
rect 686 893 688 895
rect 559 885 566 887
rect 559 883 561 885
rect 563 883 566 885
rect 515 881 518 883
rect 520 881 522 883
rect 515 879 522 881
rect 533 880 538 883
rect 515 876 520 879
rect 531 878 538 880
rect 531 876 533 878
rect 535 876 538 878
rect 531 874 538 876
rect 540 881 551 883
rect 559 881 566 883
rect 540 879 547 881
rect 549 879 551 881
rect 540 874 551 879
rect 561 876 566 881
rect 568 876 573 887
rect 575 885 584 887
rect 618 887 625 893
rect 681 888 688 893
rect 709 894 715 896
rect 709 893 717 894
rect 709 891 711 893
rect 713 891 717 893
rect 618 885 627 887
rect 575 876 586 885
rect 588 883 595 885
rect 588 881 591 883
rect 593 881 595 883
rect 588 879 595 881
rect 607 883 614 885
rect 607 881 609 883
rect 611 881 614 883
rect 607 879 614 881
rect 588 876 593 879
rect 609 876 614 879
rect 616 876 627 885
rect 629 876 634 887
rect 636 885 643 887
rect 636 883 639 885
rect 641 883 643 885
rect 636 881 643 883
rect 656 886 663 888
rect 656 884 658 886
rect 660 884 663 886
rect 656 882 663 884
rect 636 876 641 881
rect 658 875 663 882
rect 665 875 670 888
rect 672 875 677 888
rect 679 884 688 888
rect 679 875 690 884
rect 692 881 697 884
rect 692 879 699 881
rect 692 877 695 879
rect 697 877 699 879
rect 692 875 699 877
rect 709 874 717 891
rect 719 874 724 894
rect 726 874 731 894
rect 733 888 738 894
rect 733 886 740 888
rect 733 884 736 886
rect 738 884 740 886
rect 733 882 740 884
rect 733 874 738 882
rect 85 774 90 782
rect 83 772 90 774
rect 83 770 85 772
rect 87 770 90 772
rect 83 768 90 770
rect 85 762 90 768
rect 92 762 97 782
rect 99 762 104 782
rect 106 765 114 782
rect 124 779 131 781
rect 124 777 126 779
rect 128 777 131 779
rect 124 775 131 777
rect 126 772 131 775
rect 133 772 144 781
rect 135 768 144 772
rect 146 768 151 781
rect 153 768 158 781
rect 160 774 165 781
rect 182 775 187 780
rect 160 772 167 774
rect 160 770 163 772
rect 165 770 167 772
rect 160 768 167 770
rect 180 773 187 775
rect 180 771 182 773
rect 184 771 187 773
rect 180 769 187 771
rect 189 769 194 780
rect 196 771 207 780
rect 209 777 214 780
rect 230 777 235 780
rect 209 775 216 777
rect 209 773 212 775
rect 214 773 216 775
rect 209 771 216 773
rect 228 775 235 777
rect 228 773 230 775
rect 232 773 235 775
rect 228 771 235 773
rect 237 771 248 780
rect 196 769 205 771
rect 106 763 110 765
rect 112 763 114 765
rect 106 762 114 763
rect 108 760 114 762
rect 135 763 142 768
rect 198 763 205 769
rect 239 769 248 771
rect 250 769 255 780
rect 257 775 262 780
rect 272 777 283 782
rect 272 775 274 777
rect 276 775 283 777
rect 257 773 264 775
rect 272 773 283 775
rect 285 780 292 782
rect 285 778 288 780
rect 290 778 292 780
rect 285 776 292 778
rect 303 777 308 780
rect 285 773 290 776
rect 301 775 308 777
rect 301 773 303 775
rect 305 773 308 775
rect 257 771 260 773
rect 262 771 264 773
rect 257 769 264 771
rect 135 761 137 763
rect 139 761 142 763
rect 135 759 142 761
rect 198 761 201 763
rect 203 761 205 763
rect 198 759 205 761
rect 239 763 246 769
rect 301 771 308 773
rect 310 771 321 780
rect 312 769 321 771
rect 323 769 328 780
rect 330 775 335 780
rect 330 773 337 775
rect 446 774 451 781
rect 330 771 333 773
rect 335 771 337 773
rect 330 769 337 771
rect 444 772 451 774
rect 444 770 446 772
rect 448 770 451 772
rect 239 761 241 763
rect 243 761 246 763
rect 239 759 246 761
rect 312 763 319 769
rect 444 768 451 770
rect 453 768 458 781
rect 460 768 465 781
rect 467 772 478 781
rect 480 779 487 781
rect 480 777 483 779
rect 485 777 487 779
rect 480 775 487 777
rect 497 775 502 780
rect 480 772 485 775
rect 495 773 502 775
rect 467 768 476 772
rect 469 763 476 768
rect 495 771 497 773
rect 499 771 502 773
rect 495 769 502 771
rect 504 769 509 780
rect 511 771 522 780
rect 524 777 529 780
rect 539 777 550 782
rect 524 775 531 777
rect 524 773 527 775
rect 529 773 531 775
rect 539 775 541 777
rect 543 775 550 777
rect 539 773 550 775
rect 552 780 559 782
rect 552 778 555 780
rect 557 778 559 780
rect 552 776 559 778
rect 571 777 576 780
rect 552 773 557 776
rect 569 775 576 777
rect 569 773 571 775
rect 573 773 576 775
rect 524 771 531 773
rect 511 769 520 771
rect 312 761 314 763
rect 316 761 319 763
rect 312 759 319 761
rect 469 761 472 763
rect 474 761 476 763
rect 469 759 476 761
rect 513 763 520 769
rect 569 771 576 773
rect 578 771 589 780
rect 580 769 589 771
rect 591 769 596 780
rect 598 775 603 780
rect 624 775 629 780
rect 598 773 605 775
rect 598 771 601 773
rect 603 771 605 773
rect 598 769 605 771
rect 622 773 629 775
rect 622 771 624 773
rect 626 771 629 773
rect 622 769 629 771
rect 631 769 636 780
rect 638 771 649 780
rect 651 777 656 780
rect 651 775 658 777
rect 673 775 678 780
rect 651 773 654 775
rect 656 773 658 775
rect 651 771 658 773
rect 671 773 678 775
rect 671 771 673 773
rect 675 771 678 773
rect 638 769 647 771
rect 513 761 516 763
rect 518 761 520 763
rect 513 759 520 761
rect 580 763 587 769
rect 580 761 582 763
rect 584 761 587 763
rect 580 759 587 761
rect 640 763 647 769
rect 671 769 678 771
rect 680 769 685 780
rect 687 771 698 780
rect 700 777 705 780
rect 700 775 707 777
rect 700 773 703 775
rect 705 773 707 775
rect 700 771 707 773
rect 714 773 721 775
rect 714 771 716 773
rect 718 771 721 773
rect 687 769 696 771
rect 640 761 643 763
rect 645 761 647 763
rect 640 759 647 761
rect 689 763 696 769
rect 714 769 721 771
rect 689 761 692 763
rect 694 761 696 763
rect 689 759 696 761
rect 716 763 721 769
rect 723 763 728 775
rect 730 767 742 775
rect 730 765 738 767
rect 740 765 742 767
rect 730 763 742 765
rect 134 751 140 753
rect 134 749 136 751
rect 138 749 140 751
rect 134 747 140 749
rect 118 744 123 747
rect 94 742 103 744
rect 94 740 96 742
rect 98 740 103 742
rect 94 739 103 740
rect 82 736 87 739
rect 80 734 87 736
rect 80 732 82 734
rect 84 732 87 734
rect 80 730 87 732
rect 89 735 103 739
rect 105 739 113 744
rect 105 737 108 739
rect 110 737 113 739
rect 105 735 113 737
rect 115 741 123 744
rect 115 739 118 741
rect 120 739 123 741
rect 115 735 123 739
rect 125 735 130 747
rect 132 735 140 747
rect 175 745 180 749
rect 153 742 160 745
rect 153 740 155 742
rect 157 740 160 742
rect 153 738 160 740
rect 89 730 94 735
rect 155 730 160 738
rect 162 734 170 745
rect 162 732 165 734
rect 167 732 170 734
rect 162 730 170 732
rect 172 742 180 745
rect 172 740 175 742
rect 177 740 180 742
rect 172 735 180 740
rect 172 733 175 735
rect 177 733 180 735
rect 172 730 180 733
rect 182 743 189 749
rect 226 751 233 753
rect 226 749 229 751
rect 231 749 233 751
rect 182 741 185 743
rect 187 741 189 743
rect 226 743 233 749
rect 208 741 215 743
rect 182 730 191 741
rect 193 736 198 741
rect 208 739 210 741
rect 212 739 215 741
rect 208 737 215 739
rect 193 734 200 736
rect 193 732 196 734
rect 198 732 200 734
rect 210 732 215 737
rect 217 732 222 743
rect 224 741 233 743
rect 306 751 312 753
rect 306 749 308 751
rect 310 749 312 751
rect 306 747 312 749
rect 530 751 537 753
rect 530 749 532 751
rect 534 749 537 751
rect 290 744 295 747
rect 266 742 275 744
rect 224 732 235 741
rect 237 739 244 741
rect 266 740 268 742
rect 270 740 275 742
rect 266 739 275 740
rect 237 737 240 739
rect 242 737 244 739
rect 237 735 244 737
rect 254 736 259 739
rect 237 732 242 735
rect 252 734 259 736
rect 252 732 254 734
rect 256 732 259 734
rect 193 730 200 732
rect 252 730 259 732
rect 261 735 275 739
rect 277 739 285 744
rect 277 737 280 739
rect 282 737 285 739
rect 277 735 285 737
rect 287 741 295 744
rect 287 739 290 741
rect 292 739 295 741
rect 287 735 295 739
rect 297 735 302 747
rect 304 735 312 747
rect 530 743 537 749
rect 617 751 623 753
rect 617 749 619 751
rect 621 749 623 751
rect 617 747 623 749
rect 661 751 668 753
rect 661 749 664 751
rect 666 749 668 751
rect 601 744 606 747
rect 530 741 539 743
rect 519 739 526 741
rect 322 736 327 739
rect 261 730 266 735
rect 320 734 327 736
rect 320 732 322 734
rect 324 732 327 734
rect 320 730 327 732
rect 329 737 340 739
rect 329 735 336 737
rect 338 735 340 737
rect 519 737 521 739
rect 523 737 526 739
rect 519 735 526 737
rect 329 730 340 735
rect 521 732 526 735
rect 528 732 539 741
rect 541 732 546 743
rect 548 741 555 743
rect 548 739 551 741
rect 553 739 555 741
rect 577 742 586 744
rect 577 740 579 742
rect 581 740 586 742
rect 577 739 586 740
rect 548 737 555 739
rect 548 732 553 737
rect 565 736 570 739
rect 563 734 570 736
rect 563 732 565 734
rect 567 732 570 734
rect 563 730 570 732
rect 572 735 586 739
rect 588 739 596 744
rect 588 737 591 739
rect 593 737 596 739
rect 588 735 596 737
rect 598 741 606 744
rect 598 739 601 741
rect 603 739 606 741
rect 598 735 606 739
rect 608 735 613 747
rect 615 735 623 747
rect 661 743 668 749
rect 737 751 743 753
rect 737 749 739 751
rect 741 749 743 751
rect 643 741 650 743
rect 643 739 645 741
rect 647 739 650 741
rect 643 737 650 739
rect 572 730 577 735
rect 645 732 650 737
rect 652 732 657 743
rect 659 741 668 743
rect 659 732 670 741
rect 672 739 679 741
rect 737 744 743 749
rect 726 742 733 744
rect 726 741 728 742
rect 715 739 722 741
rect 672 737 675 739
rect 677 737 679 739
rect 672 735 679 737
rect 687 737 698 739
rect 687 735 689 737
rect 691 735 698 737
rect 672 732 677 735
rect 687 730 698 735
rect 700 736 705 739
rect 715 737 717 739
rect 719 737 722 739
rect 700 734 707 736
rect 700 732 703 734
rect 705 732 707 734
rect 715 733 722 737
rect 724 740 728 741
rect 730 740 733 742
rect 724 736 733 740
rect 735 743 743 744
rect 735 739 746 743
rect 735 736 743 739
rect 724 733 729 736
rect 700 730 707 732
rect 130 633 141 638
rect 81 622 89 633
rect 81 620 84 622
rect 86 620 89 622
rect 81 618 89 620
rect 91 629 99 633
rect 91 627 94 629
rect 96 627 99 629
rect 91 618 99 627
rect 101 629 109 633
rect 130 631 132 633
rect 134 631 141 633
rect 101 627 104 629
rect 106 627 109 629
rect 101 622 109 627
rect 101 620 104 622
rect 106 620 109 622
rect 101 618 109 620
rect 130 629 141 631
rect 143 636 150 638
rect 143 634 146 636
rect 148 634 150 636
rect 143 632 150 634
rect 162 633 167 636
rect 143 629 148 632
rect 160 631 167 633
rect 160 629 162 631
rect 164 629 167 631
rect 160 627 167 629
rect 169 627 180 636
rect 171 625 180 627
rect 182 625 187 636
rect 189 631 194 636
rect 515 635 522 637
rect 515 633 517 635
rect 519 633 522 635
rect 189 629 196 631
rect 189 627 192 629
rect 194 627 196 629
rect 189 625 196 627
rect 171 619 178 625
rect 205 622 213 633
rect 205 620 208 622
rect 210 620 213 622
rect 171 617 173 619
rect 175 617 178 619
rect 205 618 213 620
rect 215 629 223 633
rect 215 627 218 629
rect 220 627 223 629
rect 215 618 223 627
rect 225 629 233 633
rect 515 631 522 633
rect 225 627 228 629
rect 230 627 233 629
rect 225 622 233 627
rect 225 620 228 622
rect 230 620 233 622
rect 225 618 233 620
rect 517 628 522 631
rect 524 628 535 637
rect 526 624 535 628
rect 537 624 542 637
rect 544 624 549 637
rect 551 630 556 637
rect 551 628 558 630
rect 551 626 554 628
rect 556 626 558 628
rect 551 624 558 626
rect 575 628 582 630
rect 575 626 577 628
rect 579 626 582 628
rect 575 624 582 626
rect 171 615 178 617
rect 526 619 533 624
rect 577 620 582 624
rect 584 620 594 630
rect 596 628 604 630
rect 596 626 599 628
rect 601 626 604 628
rect 596 620 604 626
rect 606 620 615 630
rect 526 617 528 619
rect 530 617 533 619
rect 526 615 533 617
rect 586 619 592 620
rect 586 617 588 619
rect 590 617 592 619
rect 586 615 592 617
rect 608 619 615 620
rect 608 617 610 619
rect 612 617 615 619
rect 608 615 615 617
rect 647 629 656 638
rect 647 627 649 629
rect 651 627 656 629
rect 647 622 656 627
rect 647 620 649 622
rect 651 620 656 622
rect 647 618 656 620
rect 658 618 663 638
rect 665 630 670 638
rect 729 633 734 638
rect 665 628 672 630
rect 665 626 668 628
rect 670 626 672 628
rect 665 624 672 626
rect 665 618 670 624
rect 683 621 691 633
rect 693 621 698 633
rect 700 629 708 633
rect 700 627 703 629
rect 705 627 708 629
rect 700 624 708 627
rect 710 631 718 633
rect 710 629 713 631
rect 715 629 718 631
rect 710 624 718 629
rect 720 629 734 633
rect 736 636 743 638
rect 736 634 739 636
rect 741 634 743 636
rect 736 632 743 634
rect 736 629 741 632
rect 720 628 729 629
rect 720 626 725 628
rect 727 626 729 628
rect 720 624 729 626
rect 700 621 705 624
rect 683 619 689 621
rect 683 617 685 619
rect 687 617 689 619
rect 683 615 689 617
rect 134 607 140 609
rect 134 605 136 607
rect 138 605 140 607
rect 204 607 211 609
rect 134 603 140 605
rect 118 600 123 603
rect 94 598 103 600
rect 94 596 96 598
rect 98 596 103 598
rect 94 595 103 596
rect 82 592 87 595
rect 80 590 87 592
rect 80 588 82 590
rect 84 588 87 590
rect 80 586 87 588
rect 89 591 103 595
rect 105 595 113 600
rect 105 593 108 595
rect 110 593 113 595
rect 105 591 113 593
rect 115 597 123 600
rect 115 595 118 597
rect 120 595 123 597
rect 115 591 123 595
rect 125 591 130 603
rect 132 591 140 603
rect 153 600 158 606
rect 151 598 158 600
rect 151 596 153 598
rect 155 596 158 598
rect 151 594 158 596
rect 89 586 94 591
rect 153 586 158 594
rect 160 586 165 606
rect 167 604 176 606
rect 204 605 207 607
rect 209 605 211 607
rect 167 602 172 604
rect 174 602 176 604
rect 167 597 176 602
rect 204 599 211 605
rect 540 607 546 609
rect 540 605 542 607
rect 544 605 546 607
rect 617 607 624 609
rect 617 605 620 607
rect 622 605 624 607
rect 167 595 172 597
rect 174 595 176 597
rect 167 586 176 595
rect 186 597 193 599
rect 186 595 188 597
rect 190 595 193 597
rect 186 593 193 595
rect 188 588 193 593
rect 195 588 200 599
rect 202 597 211 599
rect 202 588 213 597
rect 215 595 222 597
rect 215 593 218 595
rect 220 593 222 595
rect 215 591 222 593
rect 236 592 241 595
rect 215 588 220 591
rect 234 590 241 592
rect 234 588 236 590
rect 238 588 241 590
rect 234 586 241 588
rect 243 593 254 595
rect 243 591 250 593
rect 252 591 254 593
rect 243 586 254 591
rect 540 600 546 605
rect 617 600 624 605
rect 661 607 668 609
rect 661 605 664 607
rect 666 605 668 607
rect 519 598 526 600
rect 519 596 521 598
rect 523 596 526 598
rect 519 594 526 596
rect 528 598 536 600
rect 528 596 531 598
rect 533 596 536 598
rect 528 594 536 596
rect 538 594 548 600
rect 550 598 558 600
rect 550 596 553 598
rect 555 596 558 598
rect 550 594 558 596
rect 560 598 567 600
rect 560 596 563 598
rect 565 596 567 598
rect 560 594 567 596
rect 592 598 599 600
rect 592 596 594 598
rect 596 596 599 598
rect 592 594 599 596
rect 594 587 599 594
rect 601 587 606 600
rect 608 587 613 600
rect 615 596 624 600
rect 661 599 668 605
rect 715 604 724 606
rect 715 602 717 604
rect 719 602 724 604
rect 643 597 650 599
rect 615 587 626 596
rect 628 593 633 596
rect 643 595 645 597
rect 647 595 650 597
rect 643 593 650 595
rect 628 591 635 593
rect 628 589 631 591
rect 633 589 635 591
rect 628 587 635 589
rect 645 588 650 593
rect 652 588 657 599
rect 659 597 668 599
rect 659 588 670 597
rect 672 595 679 597
rect 715 597 724 602
rect 715 595 717 597
rect 719 595 724 597
rect 672 593 675 595
rect 677 593 679 595
rect 672 591 679 593
rect 687 593 698 595
rect 687 591 689 593
rect 691 591 698 593
rect 672 588 677 591
rect 687 586 698 591
rect 700 592 705 595
rect 700 590 707 592
rect 700 588 703 590
rect 705 588 707 590
rect 700 586 707 588
rect 715 586 724 595
rect 726 586 731 606
rect 733 600 738 606
rect 733 598 740 600
rect 733 596 736 598
rect 738 596 740 598
rect 733 594 740 596
rect 733 586 738 594
rect 128 489 139 494
rect 81 478 89 489
rect 81 476 84 478
rect 86 476 89 478
rect 81 474 89 476
rect 91 485 99 489
rect 91 483 94 485
rect 96 483 99 485
rect 91 474 99 483
rect 101 485 109 489
rect 128 487 130 489
rect 132 487 139 489
rect 101 483 104 485
rect 106 483 109 485
rect 101 478 109 483
rect 101 476 104 478
rect 106 476 109 478
rect 101 474 109 476
rect 128 485 139 487
rect 141 492 148 494
rect 141 490 144 492
rect 146 490 148 492
rect 141 488 148 490
rect 205 489 210 494
rect 141 485 146 488
rect 159 477 167 489
rect 169 477 174 489
rect 176 485 184 489
rect 176 483 179 485
rect 181 483 184 485
rect 176 480 184 483
rect 186 487 194 489
rect 186 485 189 487
rect 191 485 194 487
rect 186 480 194 485
rect 196 485 210 489
rect 212 492 219 494
rect 212 490 215 492
rect 217 490 219 492
rect 212 488 219 490
rect 229 488 237 494
rect 212 485 217 488
rect 229 486 231 488
rect 233 486 237 488
rect 196 484 205 485
rect 196 482 201 484
rect 203 482 205 484
rect 229 484 237 486
rect 239 492 247 494
rect 239 490 242 492
rect 244 490 247 492
rect 239 484 247 490
rect 249 485 257 494
rect 445 489 456 494
rect 445 487 447 489
rect 449 487 456 489
rect 445 485 456 487
rect 458 492 465 494
rect 458 490 461 492
rect 463 490 465 492
rect 458 488 465 490
rect 458 485 463 488
rect 249 484 253 485
rect 196 480 205 482
rect 176 477 181 480
rect 159 475 165 477
rect 159 473 161 475
rect 163 473 165 475
rect 159 471 165 473
rect 251 483 253 484
rect 255 483 257 485
rect 251 481 257 483
rect 480 475 489 494
rect 480 473 483 475
rect 485 474 489 475
rect 491 474 496 494
rect 498 474 503 494
rect 505 474 510 494
rect 512 486 517 494
rect 581 489 586 494
rect 512 484 519 486
rect 512 482 515 484
rect 517 482 519 484
rect 512 480 519 482
rect 512 474 517 480
rect 535 477 543 489
rect 545 477 550 489
rect 552 485 560 489
rect 552 483 555 485
rect 557 483 560 485
rect 552 480 560 483
rect 562 487 570 489
rect 562 485 565 487
rect 567 485 570 487
rect 562 480 570 485
rect 572 485 586 489
rect 588 492 595 494
rect 588 490 591 492
rect 593 490 595 492
rect 588 488 595 490
rect 588 485 593 488
rect 605 487 610 492
rect 603 485 610 487
rect 572 484 581 485
rect 572 482 577 484
rect 579 482 581 484
rect 572 480 581 482
rect 603 483 605 485
rect 607 483 610 485
rect 603 481 610 483
rect 612 481 617 492
rect 619 483 630 492
rect 632 489 637 492
rect 632 487 639 489
rect 632 485 635 487
rect 637 485 639 487
rect 632 483 639 485
rect 647 487 654 491
rect 647 485 649 487
rect 651 485 654 487
rect 647 483 654 485
rect 656 488 661 491
rect 729 489 734 494
rect 656 484 665 488
rect 656 483 660 484
rect 619 481 628 483
rect 552 477 557 480
rect 535 475 541 477
rect 485 473 487 474
rect 480 471 487 473
rect 535 473 537 475
rect 539 473 541 475
rect 535 471 541 473
rect 621 475 628 481
rect 658 482 660 483
rect 662 482 665 484
rect 658 480 665 482
rect 667 480 675 488
rect 621 473 624 475
rect 626 473 628 475
rect 621 471 628 473
rect 669 475 675 480
rect 669 473 671 475
rect 673 473 675 475
rect 669 471 675 473
rect 683 477 691 489
rect 693 477 698 489
rect 700 485 708 489
rect 700 483 703 485
rect 705 483 708 485
rect 700 480 708 483
rect 710 487 718 489
rect 710 485 713 487
rect 715 485 718 487
rect 710 480 718 485
rect 720 485 734 489
rect 736 492 743 494
rect 736 490 739 492
rect 741 490 743 492
rect 736 488 743 490
rect 736 485 741 488
rect 720 484 729 485
rect 720 482 725 484
rect 727 482 729 484
rect 720 480 729 482
rect 700 477 705 480
rect 683 475 689 477
rect 683 473 685 475
rect 687 473 689 475
rect 683 471 689 473
rect 80 357 86 359
rect 40 351 45 356
rect 18 350 25 351
rect 9 346 14 350
rect 7 344 14 346
rect 7 342 9 344
rect 11 342 14 344
rect 7 340 14 342
rect 16 349 25 350
rect 16 347 20 349
rect 22 347 25 349
rect 16 340 25 347
rect 27 344 35 351
rect 27 342 30 344
rect 32 342 35 344
rect 27 340 35 342
rect 37 349 45 351
rect 37 347 40 349
rect 42 347 45 349
rect 37 345 45 347
rect 47 353 52 356
rect 47 349 55 353
rect 47 347 50 349
rect 52 347 55 349
rect 47 345 55 347
rect 37 340 42 345
rect 50 342 55 345
rect 57 351 64 353
rect 80 355 82 357
rect 84 355 86 357
rect 80 352 86 355
rect 57 349 60 351
rect 62 349 64 351
rect 57 342 64 349
rect 70 348 75 352
rect 68 346 75 348
rect 68 344 70 346
rect 72 344 75 346
rect 68 342 75 344
rect 77 349 86 352
rect 180 357 186 359
rect 140 351 145 356
rect 118 350 125 351
rect 77 342 88 349
rect 90 346 97 349
rect 109 346 114 350
rect 90 344 93 346
rect 95 344 97 346
rect 90 342 97 344
rect 107 344 114 346
rect 107 342 109 344
rect 111 342 114 344
rect 107 340 114 342
rect 116 349 125 350
rect 116 347 120 349
rect 122 347 125 349
rect 116 340 125 347
rect 127 344 135 351
rect 127 342 130 344
rect 132 342 135 344
rect 127 340 135 342
rect 137 349 145 351
rect 137 347 140 349
rect 142 347 145 349
rect 137 345 145 347
rect 147 353 152 356
rect 147 349 155 353
rect 147 347 150 349
rect 152 347 155 349
rect 147 345 155 347
rect 137 340 142 345
rect 150 342 155 345
rect 157 351 164 353
rect 180 355 182 357
rect 184 355 186 357
rect 180 352 186 355
rect 157 349 160 351
rect 162 349 164 351
rect 157 342 164 349
rect 170 348 175 352
rect 168 346 175 348
rect 168 344 170 346
rect 172 344 175 346
rect 168 342 175 344
rect 177 349 186 352
rect 280 357 286 359
rect 240 351 245 356
rect 218 350 225 351
rect 177 342 188 349
rect 190 346 197 349
rect 209 346 214 350
rect 190 344 193 346
rect 195 344 197 346
rect 190 342 197 344
rect 207 344 214 346
rect 207 342 209 344
rect 211 342 214 344
rect 207 340 214 342
rect 216 349 225 350
rect 216 347 220 349
rect 222 347 225 349
rect 216 340 225 347
rect 227 344 235 351
rect 227 342 230 344
rect 232 342 235 344
rect 227 340 235 342
rect 237 349 245 351
rect 237 347 240 349
rect 242 347 245 349
rect 237 345 245 347
rect 247 353 252 356
rect 247 349 255 353
rect 247 347 250 349
rect 252 347 255 349
rect 247 345 255 347
rect 237 340 242 345
rect 250 342 255 345
rect 257 351 264 353
rect 280 355 282 357
rect 284 355 286 357
rect 280 352 286 355
rect 257 349 260 351
rect 262 349 264 351
rect 257 342 264 349
rect 270 348 275 352
rect 268 346 275 348
rect 268 344 270 346
rect 272 344 275 346
rect 268 342 275 344
rect 277 349 286 352
rect 380 357 386 359
rect 340 351 345 356
rect 318 350 325 351
rect 277 342 288 349
rect 290 346 297 349
rect 309 346 314 350
rect 290 344 293 346
rect 295 344 297 346
rect 290 342 297 344
rect 307 344 314 346
rect 307 342 309 344
rect 311 342 314 344
rect 307 340 314 342
rect 316 349 325 350
rect 316 347 320 349
rect 322 347 325 349
rect 316 340 325 347
rect 327 344 335 351
rect 327 342 330 344
rect 332 342 335 344
rect 327 340 335 342
rect 337 349 345 351
rect 337 347 340 349
rect 342 347 345 349
rect 337 345 345 347
rect 347 353 352 356
rect 347 349 355 353
rect 347 347 350 349
rect 352 347 355 349
rect 347 345 355 347
rect 337 340 342 345
rect 350 342 355 345
rect 357 351 364 353
rect 380 355 382 357
rect 384 355 386 357
rect 380 352 386 355
rect 357 349 360 351
rect 362 349 364 351
rect 357 342 364 349
rect 370 348 375 352
rect 368 346 375 348
rect 368 344 370 346
rect 372 344 375 346
rect 368 342 375 344
rect 377 349 386 352
rect 480 357 486 359
rect 440 351 445 356
rect 418 350 425 351
rect 377 342 388 349
rect 390 346 397 349
rect 409 346 414 350
rect 390 344 393 346
rect 395 344 397 346
rect 390 342 397 344
rect 407 344 414 346
rect 407 342 409 344
rect 411 342 414 344
rect 407 340 414 342
rect 416 349 425 350
rect 416 347 420 349
rect 422 347 425 349
rect 416 340 425 347
rect 427 344 435 351
rect 427 342 430 344
rect 432 342 435 344
rect 427 340 435 342
rect 437 349 445 351
rect 437 347 440 349
rect 442 347 445 349
rect 437 345 445 347
rect 447 353 452 356
rect 447 349 455 353
rect 447 347 450 349
rect 452 347 455 349
rect 447 345 455 347
rect 437 340 442 345
rect 450 342 455 345
rect 457 351 464 353
rect 480 355 482 357
rect 484 355 486 357
rect 480 352 486 355
rect 457 349 460 351
rect 462 349 464 351
rect 457 342 464 349
rect 470 348 475 352
rect 468 346 475 348
rect 468 344 470 346
rect 472 344 475 346
rect 468 342 475 344
rect 477 349 486 352
rect 580 357 586 359
rect 540 351 545 356
rect 518 350 525 351
rect 477 342 488 349
rect 490 346 497 349
rect 509 346 514 350
rect 490 344 493 346
rect 495 344 497 346
rect 490 342 497 344
rect 507 344 514 346
rect 507 342 509 344
rect 511 342 514 344
rect 507 340 514 342
rect 516 349 525 350
rect 516 347 520 349
rect 522 347 525 349
rect 516 340 525 347
rect 527 344 535 351
rect 527 342 530 344
rect 532 342 535 344
rect 527 340 535 342
rect 537 349 545 351
rect 537 347 540 349
rect 542 347 545 349
rect 537 345 545 347
rect 547 353 552 356
rect 547 349 555 353
rect 547 347 550 349
rect 552 347 555 349
rect 547 345 555 347
rect 537 340 542 345
rect 550 342 555 345
rect 557 351 564 353
rect 580 355 582 357
rect 584 355 586 357
rect 580 352 586 355
rect 557 349 560 351
rect 562 349 564 351
rect 557 342 564 349
rect 570 348 575 352
rect 568 346 575 348
rect 568 344 570 346
rect 572 344 575 346
rect 568 342 575 344
rect 577 349 586 352
rect 680 357 686 359
rect 640 351 645 356
rect 618 350 625 351
rect 577 342 588 349
rect 590 346 597 349
rect 609 346 614 350
rect 590 344 593 346
rect 595 344 597 346
rect 590 342 597 344
rect 607 344 614 346
rect 607 342 609 344
rect 611 342 614 344
rect 607 340 614 342
rect 616 349 625 350
rect 616 347 620 349
rect 622 347 625 349
rect 616 340 625 347
rect 627 344 635 351
rect 627 342 630 344
rect 632 342 635 344
rect 627 340 635 342
rect 637 349 645 351
rect 637 347 640 349
rect 642 347 645 349
rect 637 345 645 347
rect 647 353 652 356
rect 647 349 655 353
rect 647 347 650 349
rect 652 347 655 349
rect 647 345 655 347
rect 637 340 642 345
rect 650 342 655 345
rect 657 351 664 353
rect 680 355 682 357
rect 684 355 686 357
rect 680 352 686 355
rect 657 349 660 351
rect 662 349 664 351
rect 657 342 664 349
rect 670 348 675 352
rect 668 346 675 348
rect 668 344 670 346
rect 672 344 675 346
rect 668 342 675 344
rect 677 349 686 352
rect 780 357 786 359
rect 740 351 745 356
rect 718 350 725 351
rect 677 342 688 349
rect 690 346 697 349
rect 709 346 714 350
rect 690 344 693 346
rect 695 344 697 346
rect 690 342 697 344
rect 707 344 714 346
rect 707 342 709 344
rect 711 342 714 344
rect 707 340 714 342
rect 716 349 725 350
rect 716 347 720 349
rect 722 347 725 349
rect 716 340 725 347
rect 727 344 735 351
rect 727 342 730 344
rect 732 342 735 344
rect 727 340 735 342
rect 737 349 745 351
rect 737 347 740 349
rect 742 347 745 349
rect 737 345 745 347
rect 747 353 752 356
rect 747 349 755 353
rect 747 347 750 349
rect 752 347 755 349
rect 747 345 755 347
rect 737 340 742 345
rect 750 342 755 345
rect 757 351 764 353
rect 780 355 782 357
rect 784 355 786 357
rect 780 352 786 355
rect 757 349 760 351
rect 762 349 764 351
rect 757 342 764 349
rect 770 348 775 352
rect 768 346 775 348
rect 768 344 770 346
rect 772 344 775 346
rect 768 342 775 344
rect 777 349 786 352
rect 777 342 788 349
rect 790 346 797 349
rect 790 344 793 346
rect 795 344 797 346
rect 790 342 797 344
rect 5 242 12 244
rect 5 240 7 242
rect 9 240 12 242
rect 5 237 12 240
rect 14 237 25 244
rect 16 234 25 237
rect 27 242 34 244
rect 27 240 30 242
rect 32 240 34 242
rect 27 238 34 240
rect 27 234 32 238
rect 38 237 45 244
rect 38 235 40 237
rect 42 235 45 237
rect 16 231 22 234
rect 16 229 18 231
rect 20 229 22 231
rect 38 233 45 235
rect 47 241 52 244
rect 60 241 65 246
rect 47 239 55 241
rect 47 237 50 239
rect 52 237 55 239
rect 47 233 55 237
rect 50 230 55 233
rect 57 239 65 241
rect 57 237 60 239
rect 62 237 65 239
rect 57 235 65 237
rect 67 244 75 246
rect 67 242 70 244
rect 72 242 75 244
rect 67 235 75 242
rect 77 239 86 246
rect 77 237 80 239
rect 82 237 86 239
rect 77 236 86 237
rect 88 244 95 246
rect 88 242 91 244
rect 93 242 95 244
rect 88 240 95 242
rect 105 242 112 244
rect 105 240 107 242
rect 109 240 112 242
rect 88 236 93 240
rect 105 237 112 240
rect 114 237 125 244
rect 77 235 84 236
rect 57 230 62 235
rect 16 227 22 229
rect 116 234 125 237
rect 127 242 134 244
rect 127 240 130 242
rect 132 240 134 242
rect 127 238 134 240
rect 127 234 132 238
rect 138 237 145 244
rect 138 235 140 237
rect 142 235 145 237
rect 116 231 122 234
rect 116 229 118 231
rect 120 229 122 231
rect 138 233 145 235
rect 147 241 152 244
rect 160 241 165 246
rect 147 239 155 241
rect 147 237 150 239
rect 152 237 155 239
rect 147 233 155 237
rect 150 230 155 233
rect 157 239 165 241
rect 157 237 160 239
rect 162 237 165 239
rect 157 235 165 237
rect 167 244 175 246
rect 167 242 170 244
rect 172 242 175 244
rect 167 235 175 242
rect 177 239 186 246
rect 177 237 180 239
rect 182 237 186 239
rect 177 236 186 237
rect 188 244 195 246
rect 188 242 191 244
rect 193 242 195 244
rect 188 240 195 242
rect 205 242 212 244
rect 205 240 207 242
rect 209 240 212 242
rect 188 236 193 240
rect 205 237 212 240
rect 214 237 225 244
rect 177 235 184 236
rect 157 230 162 235
rect 116 227 122 229
rect 216 234 225 237
rect 227 242 234 244
rect 227 240 230 242
rect 232 240 234 242
rect 227 238 234 240
rect 227 234 232 238
rect 238 237 245 244
rect 238 235 240 237
rect 242 235 245 237
rect 216 231 222 234
rect 216 229 218 231
rect 220 229 222 231
rect 238 233 245 235
rect 247 241 252 244
rect 260 241 265 246
rect 247 239 255 241
rect 247 237 250 239
rect 252 237 255 239
rect 247 233 255 237
rect 250 230 255 233
rect 257 239 265 241
rect 257 237 260 239
rect 262 237 265 239
rect 257 235 265 237
rect 267 244 275 246
rect 267 242 270 244
rect 272 242 275 244
rect 267 235 275 242
rect 277 239 286 246
rect 277 237 280 239
rect 282 237 286 239
rect 277 236 286 237
rect 288 244 295 246
rect 288 242 291 244
rect 293 242 295 244
rect 288 240 295 242
rect 305 242 312 244
rect 305 240 307 242
rect 309 240 312 242
rect 288 236 293 240
rect 305 237 312 240
rect 314 237 325 244
rect 277 235 284 236
rect 257 230 262 235
rect 216 227 222 229
rect 316 234 325 237
rect 327 242 334 244
rect 327 240 330 242
rect 332 240 334 242
rect 327 238 334 240
rect 327 234 332 238
rect 338 237 345 244
rect 338 235 340 237
rect 342 235 345 237
rect 316 231 322 234
rect 316 229 318 231
rect 320 229 322 231
rect 338 233 345 235
rect 347 241 352 244
rect 360 241 365 246
rect 347 239 355 241
rect 347 237 350 239
rect 352 237 355 239
rect 347 233 355 237
rect 350 230 355 233
rect 357 239 365 241
rect 357 237 360 239
rect 362 237 365 239
rect 357 235 365 237
rect 367 244 375 246
rect 367 242 370 244
rect 372 242 375 244
rect 367 235 375 242
rect 377 239 386 246
rect 377 237 380 239
rect 382 237 386 239
rect 377 236 386 237
rect 388 244 395 246
rect 388 242 391 244
rect 393 242 395 244
rect 388 240 395 242
rect 407 242 414 244
rect 407 240 409 242
rect 411 240 414 242
rect 388 236 393 240
rect 407 237 414 240
rect 416 237 427 244
rect 377 235 384 236
rect 357 230 362 235
rect 316 227 322 229
rect 418 234 427 237
rect 429 242 436 244
rect 429 240 432 242
rect 434 240 436 242
rect 429 238 436 240
rect 429 234 434 238
rect 440 237 447 244
rect 440 235 442 237
rect 444 235 447 237
rect 418 231 424 234
rect 418 229 420 231
rect 422 229 424 231
rect 440 233 447 235
rect 449 241 454 244
rect 462 241 467 246
rect 449 239 457 241
rect 449 237 452 239
rect 454 237 457 239
rect 449 233 457 237
rect 452 230 457 233
rect 459 239 467 241
rect 459 237 462 239
rect 464 237 467 239
rect 459 235 467 237
rect 469 244 477 246
rect 469 242 472 244
rect 474 242 477 244
rect 469 235 477 242
rect 479 239 488 246
rect 479 237 482 239
rect 484 237 488 239
rect 479 236 488 237
rect 490 244 497 246
rect 490 242 493 244
rect 495 242 497 244
rect 490 240 497 242
rect 507 242 514 244
rect 507 240 509 242
rect 511 240 514 242
rect 490 236 495 240
rect 507 237 514 240
rect 516 237 527 244
rect 479 235 486 236
rect 459 230 464 235
rect 418 227 424 229
rect 518 234 527 237
rect 529 242 536 244
rect 529 240 532 242
rect 534 240 536 242
rect 529 238 536 240
rect 529 234 534 238
rect 540 237 547 244
rect 540 235 542 237
rect 544 235 547 237
rect 518 231 524 234
rect 518 229 520 231
rect 522 229 524 231
rect 540 233 547 235
rect 549 241 554 244
rect 562 241 567 246
rect 549 239 557 241
rect 549 237 552 239
rect 554 237 557 239
rect 549 233 557 237
rect 552 230 557 233
rect 559 239 567 241
rect 559 237 562 239
rect 564 237 567 239
rect 559 235 567 237
rect 569 244 577 246
rect 569 242 572 244
rect 574 242 577 244
rect 569 235 577 242
rect 579 239 588 246
rect 579 237 582 239
rect 584 237 588 239
rect 579 236 588 237
rect 590 244 597 246
rect 590 242 593 244
rect 595 242 597 244
rect 590 240 597 242
rect 607 242 614 244
rect 607 240 609 242
rect 611 240 614 242
rect 590 236 595 240
rect 607 237 614 240
rect 616 237 627 244
rect 579 235 586 236
rect 559 230 564 235
rect 518 227 524 229
rect 618 234 627 237
rect 629 242 636 244
rect 629 240 632 242
rect 634 240 636 242
rect 629 238 636 240
rect 629 234 634 238
rect 640 237 647 244
rect 640 235 642 237
rect 644 235 647 237
rect 618 231 624 234
rect 618 229 620 231
rect 622 229 624 231
rect 640 233 647 235
rect 649 241 654 244
rect 662 241 667 246
rect 649 239 657 241
rect 649 237 652 239
rect 654 237 657 239
rect 649 233 657 237
rect 652 230 657 233
rect 659 239 667 241
rect 659 237 662 239
rect 664 237 667 239
rect 659 235 667 237
rect 669 244 677 246
rect 669 242 672 244
rect 674 242 677 244
rect 669 235 677 242
rect 679 239 688 246
rect 679 237 682 239
rect 684 237 688 239
rect 679 236 688 237
rect 690 244 697 246
rect 690 242 693 244
rect 695 242 697 244
rect 690 240 697 242
rect 707 242 714 244
rect 707 240 709 242
rect 711 240 714 242
rect 690 236 695 240
rect 707 237 714 240
rect 716 237 727 244
rect 679 235 686 236
rect 659 230 664 235
rect 618 227 624 229
rect 718 234 727 237
rect 729 242 736 244
rect 729 240 732 242
rect 734 240 736 242
rect 729 238 736 240
rect 729 234 734 238
rect 740 237 747 244
rect 740 235 742 237
rect 744 235 747 237
rect 718 231 724 234
rect 718 229 720 231
rect 722 229 724 231
rect 740 233 747 235
rect 749 241 754 244
rect 762 241 767 246
rect 749 239 757 241
rect 749 237 752 239
rect 754 237 757 239
rect 749 233 757 237
rect 752 230 757 233
rect 759 239 767 241
rect 759 237 762 239
rect 764 237 767 239
rect 759 235 767 237
rect 769 244 777 246
rect 769 242 772 244
rect 774 242 777 244
rect 769 235 777 242
rect 779 239 788 246
rect 779 237 782 239
rect 784 237 788 239
rect 779 236 788 237
rect 790 244 797 246
rect 790 242 793 244
rect 795 242 797 244
rect 790 240 797 242
rect 790 236 795 240
rect 779 235 786 236
rect 759 230 764 235
rect 718 227 724 229
rect 16 213 22 215
rect 16 211 18 213
rect 20 211 22 213
rect 16 208 22 211
rect 50 209 55 212
rect 16 205 25 208
rect 5 202 12 205
rect 5 200 7 202
rect 9 200 12 202
rect 5 198 12 200
rect 14 198 25 205
rect 27 204 32 208
rect 38 207 45 209
rect 38 205 40 207
rect 42 205 45 207
rect 27 202 34 204
rect 27 200 30 202
rect 32 200 34 202
rect 27 198 34 200
rect 38 198 45 205
rect 47 205 55 209
rect 47 203 50 205
rect 52 203 55 205
rect 47 201 55 203
rect 57 207 62 212
rect 57 205 65 207
rect 57 203 60 205
rect 62 203 65 205
rect 57 201 65 203
rect 47 198 52 201
rect 60 196 65 201
rect 67 200 75 207
rect 67 198 70 200
rect 72 198 75 200
rect 67 196 75 198
rect 77 206 84 207
rect 77 205 86 206
rect 77 203 80 205
rect 82 203 86 205
rect 77 196 86 203
rect 88 202 93 206
rect 116 213 122 215
rect 116 211 118 213
rect 120 211 122 213
rect 116 208 122 211
rect 150 209 155 212
rect 116 205 125 208
rect 105 202 112 205
rect 88 200 95 202
rect 88 198 91 200
rect 93 198 95 200
rect 105 200 107 202
rect 109 200 112 202
rect 105 198 112 200
rect 114 198 125 205
rect 127 204 132 208
rect 138 207 145 209
rect 138 205 140 207
rect 142 205 145 207
rect 127 202 134 204
rect 127 200 130 202
rect 132 200 134 202
rect 127 198 134 200
rect 138 198 145 205
rect 147 205 155 209
rect 147 203 150 205
rect 152 203 155 205
rect 147 201 155 203
rect 157 207 162 212
rect 157 205 165 207
rect 157 203 160 205
rect 162 203 165 205
rect 157 201 165 203
rect 147 198 152 201
rect 88 196 95 198
rect 160 196 165 201
rect 167 200 175 207
rect 167 198 170 200
rect 172 198 175 200
rect 167 196 175 198
rect 177 206 184 207
rect 177 205 186 206
rect 177 203 180 205
rect 182 203 186 205
rect 177 196 186 203
rect 188 202 193 206
rect 216 213 222 215
rect 216 211 218 213
rect 220 211 222 213
rect 216 208 222 211
rect 250 209 255 212
rect 216 205 225 208
rect 205 202 212 205
rect 188 200 195 202
rect 188 198 191 200
rect 193 198 195 200
rect 205 200 207 202
rect 209 200 212 202
rect 205 198 212 200
rect 214 198 225 205
rect 227 204 232 208
rect 238 207 245 209
rect 238 205 240 207
rect 242 205 245 207
rect 227 202 234 204
rect 227 200 230 202
rect 232 200 234 202
rect 227 198 234 200
rect 238 198 245 205
rect 247 205 255 209
rect 247 203 250 205
rect 252 203 255 205
rect 247 201 255 203
rect 257 207 262 212
rect 257 205 265 207
rect 257 203 260 205
rect 262 203 265 205
rect 257 201 265 203
rect 247 198 252 201
rect 188 196 195 198
rect 260 196 265 201
rect 267 200 275 207
rect 267 198 270 200
rect 272 198 275 200
rect 267 196 275 198
rect 277 206 284 207
rect 277 205 286 206
rect 277 203 280 205
rect 282 203 286 205
rect 277 196 286 203
rect 288 202 293 206
rect 316 213 322 215
rect 316 211 318 213
rect 320 211 322 213
rect 316 208 322 211
rect 350 209 355 212
rect 316 205 325 208
rect 305 202 312 205
rect 288 200 295 202
rect 288 198 291 200
rect 293 198 295 200
rect 305 200 307 202
rect 309 200 312 202
rect 305 198 312 200
rect 314 198 325 205
rect 327 204 332 208
rect 338 207 345 209
rect 338 205 340 207
rect 342 205 345 207
rect 327 202 334 204
rect 327 200 330 202
rect 332 200 334 202
rect 327 198 334 200
rect 338 198 345 205
rect 347 205 355 209
rect 347 203 350 205
rect 352 203 355 205
rect 347 201 355 203
rect 357 207 362 212
rect 357 205 365 207
rect 357 203 360 205
rect 362 203 365 205
rect 357 201 365 203
rect 347 198 352 201
rect 288 196 295 198
rect 360 196 365 201
rect 367 200 375 207
rect 367 198 370 200
rect 372 198 375 200
rect 367 196 375 198
rect 377 206 384 207
rect 377 205 386 206
rect 377 203 380 205
rect 382 203 386 205
rect 377 196 386 203
rect 388 202 393 206
rect 418 213 424 215
rect 418 211 420 213
rect 422 211 424 213
rect 418 208 424 211
rect 452 209 457 212
rect 418 205 427 208
rect 407 202 414 205
rect 388 200 395 202
rect 388 198 391 200
rect 393 198 395 200
rect 407 200 409 202
rect 411 200 414 202
rect 407 198 414 200
rect 416 198 427 205
rect 429 204 434 208
rect 440 207 447 209
rect 440 205 442 207
rect 444 205 447 207
rect 429 202 436 204
rect 429 200 432 202
rect 434 200 436 202
rect 429 198 436 200
rect 440 198 447 205
rect 449 205 457 209
rect 449 203 452 205
rect 454 203 457 205
rect 449 201 457 203
rect 459 207 464 212
rect 459 205 467 207
rect 459 203 462 205
rect 464 203 467 205
rect 459 201 467 203
rect 449 198 454 201
rect 388 196 395 198
rect 462 196 467 201
rect 469 200 477 207
rect 469 198 472 200
rect 474 198 477 200
rect 469 196 477 198
rect 479 206 486 207
rect 479 205 488 206
rect 479 203 482 205
rect 484 203 488 205
rect 479 196 488 203
rect 490 202 495 206
rect 518 213 524 215
rect 518 211 520 213
rect 522 211 524 213
rect 518 208 524 211
rect 552 209 557 212
rect 518 205 527 208
rect 507 202 514 205
rect 490 200 497 202
rect 490 198 493 200
rect 495 198 497 200
rect 507 200 509 202
rect 511 200 514 202
rect 507 198 514 200
rect 516 198 527 205
rect 529 204 534 208
rect 540 207 547 209
rect 540 205 542 207
rect 544 205 547 207
rect 529 202 536 204
rect 529 200 532 202
rect 534 200 536 202
rect 529 198 536 200
rect 540 198 547 205
rect 549 205 557 209
rect 549 203 552 205
rect 554 203 557 205
rect 549 201 557 203
rect 559 207 564 212
rect 559 205 567 207
rect 559 203 562 205
rect 564 203 567 205
rect 559 201 567 203
rect 549 198 554 201
rect 490 196 497 198
rect 562 196 567 201
rect 569 200 577 207
rect 569 198 572 200
rect 574 198 577 200
rect 569 196 577 198
rect 579 206 586 207
rect 579 205 588 206
rect 579 203 582 205
rect 584 203 588 205
rect 579 196 588 203
rect 590 202 595 206
rect 618 213 624 215
rect 618 211 620 213
rect 622 211 624 213
rect 618 208 624 211
rect 652 209 657 212
rect 618 205 627 208
rect 607 202 614 205
rect 590 200 597 202
rect 590 198 593 200
rect 595 198 597 200
rect 607 200 609 202
rect 611 200 614 202
rect 607 198 614 200
rect 616 198 627 205
rect 629 204 634 208
rect 640 207 647 209
rect 640 205 642 207
rect 644 205 647 207
rect 629 202 636 204
rect 629 200 632 202
rect 634 200 636 202
rect 629 198 636 200
rect 640 198 647 205
rect 649 205 657 209
rect 649 203 652 205
rect 654 203 657 205
rect 649 201 657 203
rect 659 207 664 212
rect 659 205 667 207
rect 659 203 662 205
rect 664 203 667 205
rect 659 201 667 203
rect 649 198 654 201
rect 590 196 597 198
rect 662 196 667 201
rect 669 200 677 207
rect 669 198 672 200
rect 674 198 677 200
rect 669 196 677 198
rect 679 206 686 207
rect 679 205 688 206
rect 679 203 682 205
rect 684 203 688 205
rect 679 196 688 203
rect 690 202 695 206
rect 718 213 724 215
rect 718 211 720 213
rect 722 211 724 213
rect 718 208 724 211
rect 752 209 757 212
rect 718 205 727 208
rect 707 202 714 205
rect 690 200 697 202
rect 690 198 693 200
rect 695 198 697 200
rect 707 200 709 202
rect 711 200 714 202
rect 707 198 714 200
rect 716 198 727 205
rect 729 204 734 208
rect 740 207 747 209
rect 740 205 742 207
rect 744 205 747 207
rect 729 202 736 204
rect 729 200 732 202
rect 734 200 736 202
rect 729 198 736 200
rect 740 198 747 205
rect 749 205 757 209
rect 749 203 752 205
rect 754 203 757 205
rect 749 201 757 203
rect 759 207 764 212
rect 759 205 767 207
rect 759 203 762 205
rect 764 203 767 205
rect 759 201 767 203
rect 749 198 754 201
rect 690 196 697 198
rect 762 196 767 201
rect 769 200 777 207
rect 769 198 772 200
rect 774 198 777 200
rect 769 196 777 198
rect 779 206 786 207
rect 779 205 788 206
rect 779 203 782 205
rect 784 203 788 205
rect 779 196 788 203
rect 790 202 795 206
rect 790 200 797 202
rect 790 198 793 200
rect 795 198 797 200
rect 790 196 797 198
rect 5 98 12 100
rect 5 96 7 98
rect 9 96 12 98
rect 5 93 12 96
rect 14 93 25 100
rect 16 90 25 93
rect 27 98 34 100
rect 27 96 30 98
rect 32 96 34 98
rect 27 94 34 96
rect 27 90 32 94
rect 38 93 45 100
rect 38 91 40 93
rect 42 91 45 93
rect 16 87 22 90
rect 16 85 18 87
rect 20 85 22 87
rect 38 89 45 91
rect 47 97 52 100
rect 60 97 65 102
rect 47 95 55 97
rect 47 93 50 95
rect 52 93 55 95
rect 47 89 55 93
rect 50 86 55 89
rect 57 95 65 97
rect 57 93 60 95
rect 62 93 65 95
rect 57 91 65 93
rect 67 100 75 102
rect 67 98 70 100
rect 72 98 75 100
rect 67 91 75 98
rect 77 95 86 102
rect 77 93 80 95
rect 82 93 86 95
rect 77 92 86 93
rect 88 100 95 102
rect 88 98 91 100
rect 93 98 95 100
rect 88 96 95 98
rect 105 98 112 100
rect 105 96 107 98
rect 109 96 112 98
rect 88 92 93 96
rect 105 93 112 96
rect 114 93 125 100
rect 77 91 84 92
rect 57 86 62 91
rect 16 83 22 85
rect 116 90 125 93
rect 127 98 134 100
rect 127 96 130 98
rect 132 96 134 98
rect 127 94 134 96
rect 127 90 132 94
rect 138 93 145 100
rect 138 91 140 93
rect 142 91 145 93
rect 116 87 122 90
rect 116 85 118 87
rect 120 85 122 87
rect 138 89 145 91
rect 147 97 152 100
rect 160 97 165 102
rect 147 95 155 97
rect 147 93 150 95
rect 152 93 155 95
rect 147 89 155 93
rect 150 86 155 89
rect 157 95 165 97
rect 157 93 160 95
rect 162 93 165 95
rect 157 91 165 93
rect 167 100 175 102
rect 167 98 170 100
rect 172 98 175 100
rect 167 91 175 98
rect 177 95 186 102
rect 177 93 180 95
rect 182 93 186 95
rect 177 92 186 93
rect 188 100 195 102
rect 188 98 191 100
rect 193 98 195 100
rect 188 96 195 98
rect 205 98 212 100
rect 205 96 207 98
rect 209 96 212 98
rect 188 92 193 96
rect 205 93 212 96
rect 214 93 225 100
rect 177 91 184 92
rect 157 86 162 91
rect 116 83 122 85
rect 216 90 225 93
rect 227 98 234 100
rect 227 96 230 98
rect 232 96 234 98
rect 227 94 234 96
rect 227 90 232 94
rect 238 93 245 100
rect 238 91 240 93
rect 242 91 245 93
rect 216 87 222 90
rect 216 85 218 87
rect 220 85 222 87
rect 238 89 245 91
rect 247 97 252 100
rect 260 97 265 102
rect 247 95 255 97
rect 247 93 250 95
rect 252 93 255 95
rect 247 89 255 93
rect 250 86 255 89
rect 257 95 265 97
rect 257 93 260 95
rect 262 93 265 95
rect 257 91 265 93
rect 267 100 275 102
rect 267 98 270 100
rect 272 98 275 100
rect 267 91 275 98
rect 277 95 286 102
rect 277 93 280 95
rect 282 93 286 95
rect 277 92 286 93
rect 288 100 295 102
rect 288 98 291 100
rect 293 98 295 100
rect 288 96 295 98
rect 305 98 312 100
rect 305 96 307 98
rect 309 96 312 98
rect 288 92 293 96
rect 305 93 312 96
rect 314 93 325 100
rect 277 91 284 92
rect 257 86 262 91
rect 216 83 222 85
rect 316 90 325 93
rect 327 98 334 100
rect 327 96 330 98
rect 332 96 334 98
rect 327 94 334 96
rect 327 90 332 94
rect 338 93 345 100
rect 338 91 340 93
rect 342 91 345 93
rect 316 87 322 90
rect 316 85 318 87
rect 320 85 322 87
rect 338 89 345 91
rect 347 97 352 100
rect 360 97 365 102
rect 347 95 355 97
rect 347 93 350 95
rect 352 93 355 95
rect 347 89 355 93
rect 350 86 355 89
rect 357 95 365 97
rect 357 93 360 95
rect 362 93 365 95
rect 357 91 365 93
rect 367 100 375 102
rect 367 98 370 100
rect 372 98 375 100
rect 367 91 375 98
rect 377 95 386 102
rect 377 93 380 95
rect 382 93 386 95
rect 377 92 386 93
rect 388 100 395 102
rect 388 98 391 100
rect 393 98 395 100
rect 388 96 395 98
rect 407 98 414 100
rect 407 96 409 98
rect 411 96 414 98
rect 388 92 393 96
rect 407 93 414 96
rect 416 93 427 100
rect 377 91 384 92
rect 357 86 362 91
rect 316 83 322 85
rect 418 90 427 93
rect 429 98 436 100
rect 429 96 432 98
rect 434 96 436 98
rect 429 94 436 96
rect 429 90 434 94
rect 440 93 447 100
rect 440 91 442 93
rect 444 91 447 93
rect 418 87 424 90
rect 418 85 420 87
rect 422 85 424 87
rect 440 89 447 91
rect 449 97 454 100
rect 462 97 467 102
rect 449 95 457 97
rect 449 93 452 95
rect 454 93 457 95
rect 449 89 457 93
rect 452 86 457 89
rect 459 95 467 97
rect 459 93 462 95
rect 464 93 467 95
rect 459 91 467 93
rect 469 100 477 102
rect 469 98 472 100
rect 474 98 477 100
rect 469 91 477 98
rect 479 95 488 102
rect 479 93 482 95
rect 484 93 488 95
rect 479 92 488 93
rect 490 100 497 102
rect 490 98 493 100
rect 495 98 497 100
rect 490 96 497 98
rect 507 98 514 100
rect 507 96 509 98
rect 511 96 514 98
rect 490 92 495 96
rect 507 93 514 96
rect 516 93 527 100
rect 479 91 486 92
rect 459 86 464 91
rect 418 83 424 85
rect 518 90 527 93
rect 529 98 536 100
rect 529 96 532 98
rect 534 96 536 98
rect 529 94 536 96
rect 529 90 534 94
rect 540 93 547 100
rect 540 91 542 93
rect 544 91 547 93
rect 518 87 524 90
rect 518 85 520 87
rect 522 85 524 87
rect 540 89 547 91
rect 549 97 554 100
rect 562 97 567 102
rect 549 95 557 97
rect 549 93 552 95
rect 554 93 557 95
rect 549 89 557 93
rect 552 86 557 89
rect 559 95 567 97
rect 559 93 562 95
rect 564 93 567 95
rect 559 91 567 93
rect 569 100 577 102
rect 569 98 572 100
rect 574 98 577 100
rect 569 91 577 98
rect 579 95 588 102
rect 579 93 582 95
rect 584 93 588 95
rect 579 92 588 93
rect 590 100 597 102
rect 590 98 593 100
rect 595 98 597 100
rect 590 96 597 98
rect 607 98 614 100
rect 607 96 609 98
rect 611 96 614 98
rect 590 92 595 96
rect 607 93 614 96
rect 616 93 627 100
rect 579 91 586 92
rect 559 86 564 91
rect 518 83 524 85
rect 618 90 627 93
rect 629 98 636 100
rect 629 96 632 98
rect 634 96 636 98
rect 629 94 636 96
rect 629 90 634 94
rect 640 93 647 100
rect 640 91 642 93
rect 644 91 647 93
rect 618 87 624 90
rect 618 85 620 87
rect 622 85 624 87
rect 640 89 647 91
rect 649 97 654 100
rect 662 97 667 102
rect 649 95 657 97
rect 649 93 652 95
rect 654 93 657 95
rect 649 89 657 93
rect 652 86 657 89
rect 659 95 667 97
rect 659 93 662 95
rect 664 93 667 95
rect 659 91 667 93
rect 669 100 677 102
rect 669 98 672 100
rect 674 98 677 100
rect 669 91 677 98
rect 679 95 688 102
rect 679 93 682 95
rect 684 93 688 95
rect 679 92 688 93
rect 690 100 697 102
rect 690 98 693 100
rect 695 98 697 100
rect 690 96 697 98
rect 707 98 714 100
rect 707 96 709 98
rect 711 96 714 98
rect 690 92 695 96
rect 707 93 714 96
rect 716 93 727 100
rect 679 91 686 92
rect 659 86 664 91
rect 618 83 624 85
rect 718 90 727 93
rect 729 98 736 100
rect 729 96 732 98
rect 734 96 736 98
rect 729 94 736 96
rect 729 90 734 94
rect 740 93 747 100
rect 740 91 742 93
rect 744 91 747 93
rect 718 87 724 90
rect 718 85 720 87
rect 722 85 724 87
rect 740 89 747 91
rect 749 97 754 100
rect 762 97 767 102
rect 749 95 757 97
rect 749 93 752 95
rect 754 93 757 95
rect 749 89 757 93
rect 752 86 757 89
rect 759 95 767 97
rect 759 93 762 95
rect 764 93 767 95
rect 759 91 767 93
rect 769 100 777 102
rect 769 98 772 100
rect 774 98 777 100
rect 769 91 777 98
rect 779 95 788 102
rect 779 93 782 95
rect 784 93 788 95
rect 779 92 788 93
rect 790 100 797 102
rect 790 98 793 100
rect 795 98 797 100
rect 790 96 797 98
rect 790 92 795 96
rect 779 91 786 92
rect 759 86 764 91
rect 718 83 724 85
rect 80 69 86 71
rect 40 63 45 68
rect 18 62 25 63
rect 9 58 14 62
rect 7 56 14 58
rect 7 54 9 56
rect 11 54 14 56
rect 7 52 14 54
rect 16 61 25 62
rect 16 59 20 61
rect 22 59 25 61
rect 16 52 25 59
rect 27 56 35 63
rect 27 54 30 56
rect 32 54 35 56
rect 27 52 35 54
rect 37 61 45 63
rect 37 59 40 61
rect 42 59 45 61
rect 37 57 45 59
rect 47 65 52 68
rect 47 61 55 65
rect 47 59 50 61
rect 52 59 55 61
rect 47 57 55 59
rect 37 52 42 57
rect 50 54 55 57
rect 57 63 64 65
rect 80 67 82 69
rect 84 67 86 69
rect 80 64 86 67
rect 57 61 60 63
rect 62 61 64 63
rect 57 54 64 61
rect 70 60 75 64
rect 68 58 75 60
rect 68 56 70 58
rect 72 56 75 58
rect 68 54 75 56
rect 77 61 86 64
rect 180 69 186 71
rect 140 63 145 68
rect 118 62 125 63
rect 77 54 88 61
rect 90 58 97 61
rect 109 58 114 62
rect 90 56 93 58
rect 95 56 97 58
rect 90 54 97 56
rect 107 56 114 58
rect 107 54 109 56
rect 111 54 114 56
rect 107 52 114 54
rect 116 61 125 62
rect 116 59 120 61
rect 122 59 125 61
rect 116 52 125 59
rect 127 56 135 63
rect 127 54 130 56
rect 132 54 135 56
rect 127 52 135 54
rect 137 61 145 63
rect 137 59 140 61
rect 142 59 145 61
rect 137 57 145 59
rect 147 65 152 68
rect 147 61 155 65
rect 147 59 150 61
rect 152 59 155 61
rect 147 57 155 59
rect 137 52 142 57
rect 150 54 155 57
rect 157 63 164 65
rect 180 67 182 69
rect 184 67 186 69
rect 180 64 186 67
rect 157 61 160 63
rect 162 61 164 63
rect 157 54 164 61
rect 170 60 175 64
rect 168 58 175 60
rect 168 56 170 58
rect 172 56 175 58
rect 168 54 175 56
rect 177 61 186 64
rect 280 69 286 71
rect 240 63 245 68
rect 218 62 225 63
rect 177 54 188 61
rect 190 58 197 61
rect 209 58 214 62
rect 190 56 193 58
rect 195 56 197 58
rect 190 54 197 56
rect 207 56 214 58
rect 207 54 209 56
rect 211 54 214 56
rect 207 52 214 54
rect 216 61 225 62
rect 216 59 220 61
rect 222 59 225 61
rect 216 52 225 59
rect 227 56 235 63
rect 227 54 230 56
rect 232 54 235 56
rect 227 52 235 54
rect 237 61 245 63
rect 237 59 240 61
rect 242 59 245 61
rect 237 57 245 59
rect 247 65 252 68
rect 247 61 255 65
rect 247 59 250 61
rect 252 59 255 61
rect 247 57 255 59
rect 237 52 242 57
rect 250 54 255 57
rect 257 63 264 65
rect 280 67 282 69
rect 284 67 286 69
rect 280 64 286 67
rect 257 61 260 63
rect 262 61 264 63
rect 257 54 264 61
rect 270 60 275 64
rect 268 58 275 60
rect 268 56 270 58
rect 272 56 275 58
rect 268 54 275 56
rect 277 61 286 64
rect 380 69 386 71
rect 340 63 345 68
rect 318 62 325 63
rect 277 54 288 61
rect 290 58 297 61
rect 309 58 314 62
rect 290 56 293 58
rect 295 56 297 58
rect 290 54 297 56
rect 307 56 314 58
rect 307 54 309 56
rect 311 54 314 56
rect 307 52 314 54
rect 316 61 325 62
rect 316 59 320 61
rect 322 59 325 61
rect 316 52 325 59
rect 327 56 335 63
rect 327 54 330 56
rect 332 54 335 56
rect 327 52 335 54
rect 337 61 345 63
rect 337 59 340 61
rect 342 59 345 61
rect 337 57 345 59
rect 347 65 352 68
rect 347 61 355 65
rect 347 59 350 61
rect 352 59 355 61
rect 347 57 355 59
rect 337 52 342 57
rect 350 54 355 57
rect 357 63 364 65
rect 380 67 382 69
rect 384 67 386 69
rect 380 64 386 67
rect 357 61 360 63
rect 362 61 364 63
rect 357 54 364 61
rect 370 60 375 64
rect 368 58 375 60
rect 368 56 370 58
rect 372 56 375 58
rect 368 54 375 56
rect 377 61 386 64
rect 480 69 486 71
rect 440 63 445 68
rect 418 62 425 63
rect 377 54 388 61
rect 390 58 397 61
rect 409 58 414 62
rect 390 56 393 58
rect 395 56 397 58
rect 390 54 397 56
rect 407 56 414 58
rect 407 54 409 56
rect 411 54 414 56
rect 407 52 414 54
rect 416 61 425 62
rect 416 59 420 61
rect 422 59 425 61
rect 416 52 425 59
rect 427 56 435 63
rect 427 54 430 56
rect 432 54 435 56
rect 427 52 435 54
rect 437 61 445 63
rect 437 59 440 61
rect 442 59 445 61
rect 437 57 445 59
rect 447 65 452 68
rect 447 61 455 65
rect 447 59 450 61
rect 452 59 455 61
rect 447 57 455 59
rect 437 52 442 57
rect 450 54 455 57
rect 457 63 464 65
rect 480 67 482 69
rect 484 67 486 69
rect 480 64 486 67
rect 457 61 460 63
rect 462 61 464 63
rect 457 54 464 61
rect 470 60 475 64
rect 468 58 475 60
rect 468 56 470 58
rect 472 56 475 58
rect 468 54 475 56
rect 477 61 486 64
rect 580 69 586 71
rect 540 63 545 68
rect 518 62 525 63
rect 477 54 488 61
rect 490 58 497 61
rect 509 58 514 62
rect 490 56 493 58
rect 495 56 497 58
rect 490 54 497 56
rect 507 56 514 58
rect 507 54 509 56
rect 511 54 514 56
rect 507 52 514 54
rect 516 61 525 62
rect 516 59 520 61
rect 522 59 525 61
rect 516 52 525 59
rect 527 56 535 63
rect 527 54 530 56
rect 532 54 535 56
rect 527 52 535 54
rect 537 61 545 63
rect 537 59 540 61
rect 542 59 545 61
rect 537 57 545 59
rect 547 65 552 68
rect 547 61 555 65
rect 547 59 550 61
rect 552 59 555 61
rect 547 57 555 59
rect 537 52 542 57
rect 550 54 555 57
rect 557 63 564 65
rect 580 67 582 69
rect 584 67 586 69
rect 580 64 586 67
rect 557 61 560 63
rect 562 61 564 63
rect 557 54 564 61
rect 570 60 575 64
rect 568 58 575 60
rect 568 56 570 58
rect 572 56 575 58
rect 568 54 575 56
rect 577 61 586 64
rect 680 69 686 71
rect 640 63 645 68
rect 618 62 625 63
rect 577 54 588 61
rect 590 58 597 61
rect 609 58 614 62
rect 590 56 593 58
rect 595 56 597 58
rect 590 54 597 56
rect 607 56 614 58
rect 607 54 609 56
rect 611 54 614 56
rect 607 52 614 54
rect 616 61 625 62
rect 616 59 620 61
rect 622 59 625 61
rect 616 52 625 59
rect 627 56 635 63
rect 627 54 630 56
rect 632 54 635 56
rect 627 52 635 54
rect 637 61 645 63
rect 637 59 640 61
rect 642 59 645 61
rect 637 57 645 59
rect 647 65 652 68
rect 647 61 655 65
rect 647 59 650 61
rect 652 59 655 61
rect 647 57 655 59
rect 637 52 642 57
rect 650 54 655 57
rect 657 63 664 65
rect 680 67 682 69
rect 684 67 686 69
rect 680 64 686 67
rect 657 61 660 63
rect 662 61 664 63
rect 657 54 664 61
rect 670 60 675 64
rect 668 58 675 60
rect 668 56 670 58
rect 672 56 675 58
rect 668 54 675 56
rect 677 61 686 64
rect 780 69 786 71
rect 740 63 745 68
rect 718 62 725 63
rect 677 54 688 61
rect 690 58 697 61
rect 709 58 714 62
rect 690 56 693 58
rect 695 56 697 58
rect 690 54 697 56
rect 707 56 714 58
rect 707 54 709 56
rect 711 54 714 56
rect 707 52 714 54
rect 716 61 725 62
rect 716 59 720 61
rect 722 59 725 61
rect 716 52 725 59
rect 727 56 735 63
rect 727 54 730 56
rect 732 54 735 56
rect 727 52 735 54
rect 737 61 745 63
rect 737 59 740 61
rect 742 59 745 61
rect 737 57 745 59
rect 747 65 752 68
rect 747 61 755 65
rect 747 59 750 61
rect 752 59 755 61
rect 747 57 755 59
rect 737 52 742 57
rect 750 54 755 57
rect 757 63 764 65
rect 780 67 782 69
rect 784 67 786 69
rect 780 64 786 67
rect 757 61 760 63
rect 762 61 764 63
rect 757 54 764 61
rect 770 60 775 64
rect 768 58 775 60
rect 768 56 770 58
rect 772 56 775 58
rect 768 54 775 56
rect 777 61 786 64
rect 777 54 788 61
rect 790 58 797 61
rect 790 56 793 58
rect 795 56 797 58
rect 790 54 797 56
rect -10 -72 -3 -70
rect -10 -74 -8 -72
rect -6 -74 -3 -72
rect -10 -76 -3 -74
rect -8 -80 -3 -76
rect -1 -77 8 -70
rect -1 -79 3 -77
rect 5 -79 8 -77
rect -1 -80 8 -79
rect 1 -81 8 -80
rect 10 -72 18 -70
rect 10 -74 13 -72
rect 15 -74 18 -72
rect 10 -81 18 -74
rect 20 -75 25 -70
rect 96 -72 103 -70
rect 33 -75 38 -72
rect 20 -77 28 -75
rect 20 -79 23 -77
rect 25 -79 28 -77
rect 20 -81 28 -79
rect 23 -86 28 -81
rect 30 -77 38 -75
rect 30 -79 33 -77
rect 35 -79 38 -77
rect 30 -83 38 -79
rect 40 -79 47 -72
rect 51 -74 58 -72
rect 51 -76 53 -74
rect 55 -76 58 -74
rect 51 -78 58 -76
rect 40 -81 43 -79
rect 45 -81 47 -79
rect 40 -83 47 -81
rect 53 -82 58 -78
rect 60 -79 71 -72
rect 73 -74 80 -72
rect 73 -76 76 -74
rect 78 -76 80 -74
rect 96 -74 98 -72
rect 100 -74 103 -72
rect 96 -76 103 -74
rect 73 -79 80 -76
rect 60 -82 69 -79
rect 30 -86 35 -83
rect 63 -85 69 -82
rect 63 -87 65 -85
rect 67 -87 69 -85
rect 63 -89 69 -87
rect 98 -80 103 -76
rect 105 -77 114 -70
rect 105 -79 109 -77
rect 111 -79 114 -77
rect 105 -80 114 -79
rect 107 -81 114 -80
rect 116 -72 124 -70
rect 116 -74 119 -72
rect 121 -74 124 -72
rect 116 -81 124 -74
rect 126 -75 131 -70
rect 202 -72 209 -70
rect 139 -75 144 -72
rect 126 -77 134 -75
rect 126 -79 129 -77
rect 131 -79 134 -77
rect 126 -81 134 -79
rect 129 -86 134 -81
rect 136 -77 144 -75
rect 136 -79 139 -77
rect 141 -79 144 -77
rect 136 -83 144 -79
rect 146 -79 153 -72
rect 157 -74 164 -72
rect 157 -76 159 -74
rect 161 -76 164 -74
rect 157 -78 164 -76
rect 146 -81 149 -79
rect 151 -81 153 -79
rect 146 -83 153 -81
rect 159 -82 164 -78
rect 166 -79 177 -72
rect 179 -74 186 -72
rect 179 -76 182 -74
rect 184 -76 186 -74
rect 202 -74 204 -72
rect 206 -74 209 -72
rect 202 -76 209 -74
rect 179 -79 186 -76
rect 166 -82 175 -79
rect 136 -86 141 -83
rect 169 -85 175 -82
rect 169 -87 171 -85
rect 173 -87 175 -85
rect 169 -89 175 -87
rect 204 -80 209 -76
rect 211 -77 220 -70
rect 211 -79 215 -77
rect 217 -79 220 -77
rect 211 -80 220 -79
rect 213 -81 220 -80
rect 222 -72 230 -70
rect 222 -74 225 -72
rect 227 -74 230 -72
rect 222 -81 230 -74
rect 232 -75 237 -70
rect 308 -72 315 -70
rect 245 -75 250 -72
rect 232 -77 240 -75
rect 232 -79 235 -77
rect 237 -79 240 -77
rect 232 -81 240 -79
rect 235 -86 240 -81
rect 242 -77 250 -75
rect 242 -79 245 -77
rect 247 -79 250 -77
rect 242 -83 250 -79
rect 252 -79 259 -72
rect 263 -74 270 -72
rect 263 -76 265 -74
rect 267 -76 270 -74
rect 263 -78 270 -76
rect 252 -81 255 -79
rect 257 -81 259 -79
rect 252 -83 259 -81
rect 265 -82 270 -78
rect 272 -79 283 -72
rect 285 -74 292 -72
rect 285 -76 288 -74
rect 290 -76 292 -74
rect 308 -74 310 -72
rect 312 -74 315 -72
rect 308 -76 315 -74
rect 285 -79 292 -76
rect 272 -82 281 -79
rect 242 -86 247 -83
rect 275 -85 281 -82
rect 275 -87 277 -85
rect 279 -87 281 -85
rect 275 -89 281 -87
rect 310 -80 315 -76
rect 317 -77 326 -70
rect 317 -79 321 -77
rect 323 -79 326 -77
rect 317 -80 326 -79
rect 319 -81 326 -80
rect 328 -72 336 -70
rect 328 -74 331 -72
rect 333 -74 336 -72
rect 328 -81 336 -74
rect 338 -75 343 -70
rect 414 -72 421 -70
rect 351 -75 356 -72
rect 338 -77 346 -75
rect 338 -79 341 -77
rect 343 -79 346 -77
rect 338 -81 346 -79
rect 341 -86 346 -81
rect 348 -77 356 -75
rect 348 -79 351 -77
rect 353 -79 356 -77
rect 348 -83 356 -79
rect 358 -79 365 -72
rect 369 -74 376 -72
rect 369 -76 371 -74
rect 373 -76 376 -74
rect 369 -78 376 -76
rect 358 -81 361 -79
rect 363 -81 365 -79
rect 358 -83 365 -81
rect 371 -82 376 -78
rect 378 -79 389 -72
rect 391 -74 398 -72
rect 391 -76 394 -74
rect 396 -76 398 -74
rect 414 -74 416 -72
rect 418 -74 421 -72
rect 414 -76 421 -74
rect 391 -79 398 -76
rect 378 -82 387 -79
rect 348 -86 353 -83
rect 381 -85 387 -82
rect 381 -87 383 -85
rect 385 -87 387 -85
rect 381 -89 387 -87
rect 416 -80 421 -76
rect 423 -77 432 -70
rect 423 -79 427 -77
rect 429 -79 432 -77
rect 423 -80 432 -79
rect 425 -81 432 -80
rect 434 -72 442 -70
rect 434 -74 437 -72
rect 439 -74 442 -72
rect 434 -81 442 -74
rect 444 -75 449 -70
rect 520 -72 527 -70
rect 457 -75 462 -72
rect 444 -77 452 -75
rect 444 -79 447 -77
rect 449 -79 452 -77
rect 444 -81 452 -79
rect 447 -86 452 -81
rect 454 -77 462 -75
rect 454 -79 457 -77
rect 459 -79 462 -77
rect 454 -83 462 -79
rect 464 -79 471 -72
rect 475 -74 482 -72
rect 475 -76 477 -74
rect 479 -76 482 -74
rect 475 -78 482 -76
rect 464 -81 467 -79
rect 469 -81 471 -79
rect 464 -83 471 -81
rect 477 -82 482 -78
rect 484 -79 495 -72
rect 497 -74 504 -72
rect 497 -76 500 -74
rect 502 -76 504 -74
rect 520 -74 522 -72
rect 524 -74 527 -72
rect 520 -76 527 -74
rect 497 -79 504 -76
rect 484 -82 493 -79
rect 454 -86 459 -83
rect 487 -85 493 -82
rect 487 -87 489 -85
rect 491 -87 493 -85
rect 487 -89 493 -87
rect 522 -80 527 -76
rect 529 -77 538 -70
rect 529 -79 533 -77
rect 535 -79 538 -77
rect 529 -80 538 -79
rect 531 -81 538 -80
rect 540 -72 548 -70
rect 540 -74 543 -72
rect 545 -74 548 -72
rect 540 -81 548 -74
rect 550 -75 555 -70
rect 626 -72 633 -70
rect 563 -75 568 -72
rect 550 -77 558 -75
rect 550 -79 553 -77
rect 555 -79 558 -77
rect 550 -81 558 -79
rect 553 -86 558 -81
rect 560 -77 568 -75
rect 560 -79 563 -77
rect 565 -79 568 -77
rect 560 -83 568 -79
rect 570 -79 577 -72
rect 581 -74 588 -72
rect 581 -76 583 -74
rect 585 -76 588 -74
rect 581 -78 588 -76
rect 570 -81 573 -79
rect 575 -81 577 -79
rect 570 -83 577 -81
rect 583 -82 588 -78
rect 590 -79 601 -72
rect 603 -74 610 -72
rect 603 -76 606 -74
rect 608 -76 610 -74
rect 626 -74 628 -72
rect 630 -74 633 -72
rect 626 -76 633 -74
rect 603 -79 610 -76
rect 590 -82 599 -79
rect 560 -86 565 -83
rect 593 -85 599 -82
rect 593 -87 595 -85
rect 597 -87 599 -85
rect 593 -89 599 -87
rect 628 -80 633 -76
rect 635 -77 644 -70
rect 635 -79 639 -77
rect 641 -79 644 -77
rect 635 -80 644 -79
rect 637 -81 644 -80
rect 646 -72 654 -70
rect 646 -74 649 -72
rect 651 -74 654 -72
rect 646 -81 654 -74
rect 656 -75 661 -70
rect 732 -72 739 -70
rect 669 -75 674 -72
rect 656 -77 664 -75
rect 656 -79 659 -77
rect 661 -79 664 -77
rect 656 -81 664 -79
rect 659 -86 664 -81
rect 666 -77 674 -75
rect 666 -79 669 -77
rect 671 -79 674 -77
rect 666 -83 674 -79
rect 676 -79 683 -72
rect 687 -74 694 -72
rect 687 -76 689 -74
rect 691 -76 694 -74
rect 687 -78 694 -76
rect 676 -81 679 -79
rect 681 -81 683 -79
rect 676 -83 683 -81
rect 689 -82 694 -78
rect 696 -79 707 -72
rect 709 -74 716 -72
rect 709 -76 712 -74
rect 714 -76 716 -74
rect 732 -74 734 -72
rect 736 -74 739 -72
rect 732 -76 739 -74
rect 709 -79 716 -76
rect 696 -82 705 -79
rect 666 -86 671 -83
rect 699 -85 705 -82
rect 699 -87 701 -85
rect 703 -87 705 -85
rect 699 -89 705 -87
rect 734 -80 739 -76
rect 741 -77 750 -70
rect 741 -79 745 -77
rect 747 -79 750 -77
rect 741 -80 750 -79
rect 743 -81 750 -80
rect 752 -72 760 -70
rect 752 -74 755 -72
rect 757 -74 760 -72
rect 752 -81 760 -74
rect 762 -75 767 -70
rect 838 -72 845 -70
rect 775 -75 780 -72
rect 762 -77 770 -75
rect 762 -79 765 -77
rect 767 -79 770 -77
rect 762 -81 770 -79
rect 765 -86 770 -81
rect 772 -77 780 -75
rect 772 -79 775 -77
rect 777 -79 780 -77
rect 772 -83 780 -79
rect 782 -79 789 -72
rect 793 -74 800 -72
rect 793 -76 795 -74
rect 797 -76 800 -74
rect 793 -78 800 -76
rect 782 -81 785 -79
rect 787 -81 789 -79
rect 782 -83 789 -81
rect 795 -82 800 -78
rect 802 -79 813 -72
rect 815 -74 822 -72
rect 815 -76 818 -74
rect 820 -76 822 -74
rect 838 -74 840 -72
rect 842 -74 845 -72
rect 838 -76 845 -74
rect 815 -79 822 -76
rect 802 -82 811 -79
rect 772 -86 777 -83
rect 805 -85 811 -82
rect 805 -87 807 -85
rect 809 -87 811 -85
rect 805 -89 811 -87
rect 840 -80 845 -76
rect 847 -77 856 -70
rect 847 -79 851 -77
rect 853 -79 856 -77
rect 847 -80 856 -79
rect 849 -81 856 -80
rect 858 -72 866 -70
rect 858 -74 861 -72
rect 863 -74 866 -72
rect 858 -81 866 -74
rect 868 -75 873 -70
rect 881 -75 886 -72
rect 868 -77 876 -75
rect 868 -79 871 -77
rect 873 -79 876 -77
rect 868 -81 876 -79
rect 871 -86 876 -81
rect 878 -77 886 -75
rect 878 -79 881 -77
rect 883 -79 886 -77
rect 878 -83 886 -79
rect 888 -79 895 -72
rect 899 -74 906 -72
rect 899 -76 901 -74
rect 903 -76 906 -74
rect 899 -78 906 -76
rect 888 -81 891 -79
rect 893 -81 895 -79
rect 888 -83 895 -81
rect 901 -82 906 -78
rect 908 -79 919 -72
rect 921 -74 928 -72
rect 921 -76 924 -74
rect 926 -76 928 -74
rect 921 -79 928 -76
rect 908 -82 917 -79
rect 878 -86 883 -83
rect 911 -85 917 -82
rect 911 -87 913 -85
rect 915 -87 917 -85
rect 911 -89 917 -87
<< pdif >>
rect 88 1147 95 1149
rect 88 1145 90 1147
rect 92 1145 95 1147
rect 88 1143 95 1145
rect 90 1122 95 1143
rect 97 1133 111 1149
rect 97 1131 100 1133
rect 102 1131 111 1133
rect 113 1147 121 1149
rect 113 1145 116 1147
rect 118 1145 121 1147
rect 113 1140 121 1145
rect 113 1138 116 1140
rect 118 1138 121 1140
rect 113 1131 121 1138
rect 123 1140 131 1149
rect 123 1138 126 1140
rect 128 1138 131 1140
rect 123 1131 131 1138
rect 97 1126 109 1131
rect 97 1124 100 1126
rect 102 1124 109 1126
rect 97 1122 109 1124
rect 126 1122 131 1131
rect 133 1134 138 1149
rect 153 1142 158 1150
rect 151 1140 158 1142
rect 151 1138 153 1140
rect 155 1138 158 1140
rect 133 1132 140 1134
rect 133 1130 136 1132
rect 138 1130 140 1132
rect 133 1128 140 1130
rect 151 1133 158 1138
rect 151 1131 153 1133
rect 155 1131 158 1133
rect 151 1129 158 1131
rect 133 1122 138 1128
rect 153 1122 158 1129
rect 160 1122 165 1150
rect 167 1133 176 1150
rect 184 1147 191 1149
rect 184 1145 186 1147
rect 188 1145 191 1147
rect 184 1140 191 1145
rect 184 1138 186 1140
rect 188 1138 191 1140
rect 184 1136 191 1138
rect 167 1131 172 1133
rect 174 1131 176 1133
rect 186 1131 191 1136
rect 193 1142 199 1149
rect 236 1147 243 1149
rect 236 1145 238 1147
rect 240 1145 243 1147
rect 236 1143 243 1145
rect 193 1135 201 1142
rect 193 1133 196 1135
rect 198 1133 201 1135
rect 193 1131 201 1133
rect 167 1126 176 1131
rect 195 1129 201 1131
rect 203 1140 211 1142
rect 203 1138 206 1140
rect 208 1138 211 1140
rect 203 1133 211 1138
rect 203 1131 206 1133
rect 208 1131 211 1133
rect 203 1129 211 1131
rect 213 1133 220 1142
rect 213 1131 216 1133
rect 218 1131 220 1133
rect 213 1129 220 1131
rect 167 1124 172 1126
rect 174 1124 176 1126
rect 167 1122 176 1124
rect 238 1122 243 1143
rect 245 1133 259 1149
rect 245 1131 248 1133
rect 250 1131 259 1133
rect 261 1147 269 1149
rect 261 1145 264 1147
rect 266 1145 269 1147
rect 261 1140 269 1145
rect 261 1138 264 1140
rect 266 1138 269 1140
rect 261 1131 269 1138
rect 271 1140 279 1149
rect 271 1138 274 1140
rect 276 1138 279 1140
rect 271 1131 279 1138
rect 245 1126 257 1131
rect 245 1124 248 1126
rect 250 1124 257 1126
rect 245 1122 257 1124
rect 274 1122 279 1131
rect 281 1134 286 1149
rect 358 1148 365 1150
rect 358 1146 360 1148
rect 362 1146 365 1148
rect 281 1132 288 1134
rect 281 1130 284 1132
rect 286 1130 288 1132
rect 281 1128 288 1130
rect 298 1130 305 1143
rect 298 1128 300 1130
rect 302 1128 305 1130
rect 281 1122 286 1128
rect 298 1126 305 1128
rect 307 1140 315 1143
rect 307 1138 310 1140
rect 312 1138 315 1140
rect 307 1133 315 1138
rect 307 1131 310 1133
rect 312 1131 315 1133
rect 307 1126 315 1131
rect 317 1130 325 1143
rect 317 1128 320 1130
rect 322 1128 325 1130
rect 317 1126 325 1128
rect 327 1140 335 1143
rect 327 1138 330 1140
rect 332 1138 335 1140
rect 327 1133 335 1138
rect 327 1131 330 1133
rect 332 1131 335 1133
rect 327 1126 335 1131
rect 337 1126 345 1143
rect 358 1141 365 1146
rect 358 1139 360 1141
rect 362 1139 365 1141
rect 358 1137 365 1139
rect 360 1132 365 1137
rect 367 1133 376 1150
rect 367 1132 371 1133
rect 369 1131 371 1132
rect 373 1131 376 1133
rect 369 1129 376 1131
rect 566 1134 574 1147
rect 566 1132 569 1134
rect 571 1132 574 1134
rect 566 1127 574 1132
rect 339 1123 345 1126
rect 566 1125 569 1127
rect 571 1125 574 1127
rect 339 1121 341 1123
rect 343 1121 345 1123
rect 339 1119 345 1121
rect 566 1123 574 1125
rect 576 1141 584 1147
rect 576 1139 579 1141
rect 581 1139 584 1141
rect 576 1131 584 1139
rect 586 1142 594 1147
rect 612 1147 619 1149
rect 612 1145 614 1147
rect 616 1145 619 1147
rect 612 1143 619 1145
rect 586 1140 589 1142
rect 591 1140 594 1142
rect 586 1135 594 1140
rect 586 1133 589 1135
rect 591 1133 594 1135
rect 586 1131 594 1133
rect 576 1123 581 1131
rect 614 1122 619 1143
rect 621 1133 635 1149
rect 621 1131 624 1133
rect 626 1131 635 1133
rect 637 1147 645 1149
rect 637 1145 640 1147
rect 642 1145 645 1147
rect 637 1140 645 1145
rect 637 1138 640 1140
rect 642 1138 645 1140
rect 637 1131 645 1138
rect 647 1140 655 1149
rect 647 1138 650 1140
rect 652 1138 655 1140
rect 647 1131 655 1138
rect 621 1126 633 1131
rect 621 1124 624 1126
rect 626 1124 633 1126
rect 621 1122 633 1124
rect 650 1122 655 1131
rect 657 1134 662 1149
rect 675 1148 682 1150
rect 675 1146 677 1148
rect 679 1146 682 1148
rect 675 1141 682 1146
rect 675 1139 677 1141
rect 679 1139 682 1141
rect 675 1137 682 1139
rect 657 1132 664 1134
rect 677 1132 682 1137
rect 684 1133 693 1150
rect 684 1132 688 1133
rect 657 1130 660 1132
rect 662 1130 664 1132
rect 657 1128 664 1130
rect 657 1122 662 1128
rect 686 1131 688 1132
rect 690 1131 693 1133
rect 686 1129 693 1131
rect 703 1133 710 1149
rect 703 1131 705 1133
rect 707 1131 710 1133
rect 703 1126 710 1131
rect 703 1124 705 1126
rect 707 1124 710 1126
rect 703 1122 710 1124
rect 712 1122 717 1149
rect 719 1147 727 1149
rect 719 1145 722 1147
rect 724 1145 727 1147
rect 719 1140 727 1145
rect 719 1138 722 1140
rect 724 1138 727 1140
rect 719 1122 727 1138
rect 729 1122 734 1149
rect 736 1133 743 1149
rect 736 1131 739 1133
rect 741 1131 743 1133
rect 736 1126 743 1131
rect 736 1124 739 1126
rect 741 1124 743 1126
rect 736 1122 743 1124
rect 80 1108 87 1110
rect 80 1106 82 1108
rect 84 1106 87 1108
rect 80 1101 87 1106
rect 80 1099 82 1101
rect 84 1099 87 1101
rect 80 1086 87 1099
rect 89 1101 97 1110
rect 89 1099 92 1101
rect 94 1099 97 1101
rect 89 1094 97 1099
rect 89 1092 92 1094
rect 94 1092 97 1094
rect 89 1086 97 1092
rect 99 1108 107 1110
rect 99 1106 102 1108
rect 104 1106 107 1108
rect 219 1111 225 1113
rect 219 1109 221 1111
rect 223 1109 225 1111
rect 99 1101 107 1106
rect 99 1099 102 1101
rect 104 1099 107 1101
rect 127 1101 134 1103
rect 155 1101 161 1103
rect 127 1100 129 1101
rect 99 1086 107 1099
rect 118 1095 123 1100
rect 116 1093 123 1095
rect 116 1091 118 1093
rect 120 1091 123 1093
rect 116 1086 123 1091
rect 116 1084 118 1086
rect 120 1084 123 1086
rect 116 1082 123 1084
rect 125 1099 129 1100
rect 131 1099 134 1101
rect 125 1082 134 1099
rect 146 1096 151 1101
rect 144 1094 151 1096
rect 144 1092 146 1094
rect 148 1092 151 1094
rect 144 1087 151 1092
rect 144 1085 146 1087
rect 148 1085 151 1087
rect 144 1083 151 1085
rect 153 1099 161 1101
rect 153 1097 156 1099
rect 158 1097 161 1099
rect 153 1090 161 1097
rect 163 1101 171 1103
rect 163 1099 166 1101
rect 168 1099 171 1101
rect 163 1094 171 1099
rect 163 1092 166 1094
rect 168 1092 171 1094
rect 163 1090 171 1092
rect 173 1101 180 1103
rect 219 1102 225 1109
rect 258 1111 265 1113
rect 258 1109 261 1111
rect 263 1109 265 1111
rect 258 1108 265 1109
rect 173 1099 176 1101
rect 178 1099 180 1101
rect 173 1090 180 1099
rect 190 1097 195 1102
rect 188 1095 195 1097
rect 188 1093 190 1095
rect 192 1093 195 1095
rect 153 1083 159 1090
rect 188 1088 195 1093
rect 188 1086 190 1088
rect 192 1086 195 1088
rect 188 1084 195 1086
rect 197 1100 205 1102
rect 197 1098 200 1100
rect 202 1098 205 1100
rect 197 1089 205 1098
rect 207 1100 215 1102
rect 207 1098 210 1100
rect 212 1098 215 1100
rect 207 1093 215 1098
rect 207 1091 210 1093
rect 212 1091 215 1093
rect 207 1089 215 1091
rect 217 1101 225 1102
rect 217 1089 227 1101
rect 197 1084 203 1089
rect 222 1088 227 1089
rect 229 1099 236 1101
rect 229 1097 232 1099
rect 234 1097 236 1099
rect 229 1092 236 1097
rect 229 1090 232 1092
rect 234 1090 236 1092
rect 229 1088 236 1090
rect 258 1083 267 1108
rect 269 1083 274 1108
rect 276 1083 281 1108
rect 283 1083 288 1108
rect 290 1101 295 1108
rect 648 1108 656 1110
rect 571 1101 578 1103
rect 290 1093 298 1101
rect 290 1091 293 1093
rect 295 1091 298 1093
rect 290 1083 298 1091
rect 300 1083 305 1101
rect 307 1083 312 1101
rect 314 1083 319 1101
rect 321 1099 328 1101
rect 321 1097 324 1099
rect 326 1097 328 1099
rect 321 1092 328 1097
rect 321 1090 324 1092
rect 326 1090 328 1092
rect 321 1083 328 1090
rect 571 1099 574 1101
rect 576 1100 578 1101
rect 648 1106 651 1108
rect 653 1106 656 1108
rect 612 1101 618 1103
rect 576 1099 580 1100
rect 571 1082 580 1099
rect 582 1095 587 1100
rect 603 1096 608 1101
rect 582 1093 589 1095
rect 582 1091 585 1093
rect 587 1091 589 1093
rect 582 1086 589 1091
rect 582 1084 585 1086
rect 587 1084 589 1086
rect 582 1082 589 1084
rect 601 1094 608 1096
rect 601 1092 603 1094
rect 605 1092 608 1094
rect 601 1087 608 1092
rect 601 1085 603 1087
rect 605 1085 608 1087
rect 601 1083 608 1085
rect 610 1099 618 1101
rect 610 1097 613 1099
rect 615 1097 618 1099
rect 610 1090 618 1097
rect 620 1101 628 1103
rect 620 1099 623 1101
rect 625 1099 628 1101
rect 620 1094 628 1099
rect 620 1092 623 1094
rect 625 1092 628 1094
rect 620 1090 628 1092
rect 630 1101 637 1103
rect 630 1099 633 1101
rect 635 1099 637 1101
rect 630 1090 637 1099
rect 648 1101 656 1106
rect 648 1099 651 1101
rect 653 1099 656 1101
rect 610 1083 616 1090
rect 648 1086 656 1099
rect 658 1101 666 1110
rect 658 1099 661 1101
rect 663 1099 666 1101
rect 658 1094 666 1099
rect 658 1092 661 1094
rect 663 1092 666 1094
rect 658 1086 666 1092
rect 668 1108 675 1110
rect 668 1106 671 1108
rect 673 1106 675 1108
rect 668 1101 675 1106
rect 685 1104 690 1110
rect 668 1099 671 1101
rect 673 1099 675 1101
rect 668 1086 675 1099
rect 683 1102 690 1104
rect 683 1100 685 1102
rect 687 1100 690 1102
rect 683 1098 690 1100
rect 685 1083 690 1098
rect 692 1101 697 1110
rect 714 1108 726 1110
rect 714 1106 721 1108
rect 723 1106 726 1108
rect 714 1101 726 1106
rect 692 1094 700 1101
rect 692 1092 695 1094
rect 697 1092 700 1094
rect 692 1083 700 1092
rect 702 1094 710 1101
rect 702 1092 705 1094
rect 707 1092 710 1094
rect 702 1087 710 1092
rect 702 1085 705 1087
rect 707 1085 710 1087
rect 702 1083 710 1085
rect 712 1099 721 1101
rect 723 1099 726 1101
rect 712 1083 726 1099
rect 728 1089 733 1110
rect 728 1087 735 1089
rect 728 1085 731 1087
rect 733 1085 735 1087
rect 728 1083 735 1085
rect 88 1003 95 1005
rect 88 1001 90 1003
rect 92 1001 95 1003
rect 88 999 95 1001
rect 90 978 95 999
rect 97 989 111 1005
rect 97 987 100 989
rect 102 987 111 989
rect 113 1003 121 1005
rect 113 1001 116 1003
rect 118 1001 121 1003
rect 113 996 121 1001
rect 113 994 116 996
rect 118 994 121 996
rect 113 987 121 994
rect 123 996 131 1005
rect 123 994 126 996
rect 128 994 131 996
rect 123 987 131 994
rect 97 982 109 987
rect 97 980 100 982
rect 102 980 109 982
rect 97 978 109 980
rect 126 978 131 987
rect 133 990 138 1005
rect 133 988 140 990
rect 133 986 136 988
rect 138 986 140 988
rect 133 984 140 986
rect 148 989 155 1002
rect 148 987 150 989
rect 152 987 155 989
rect 133 978 138 984
rect 148 982 155 987
rect 148 980 150 982
rect 152 980 155 982
rect 148 978 155 980
rect 157 996 165 1002
rect 157 994 160 996
rect 162 994 165 996
rect 157 989 165 994
rect 157 987 160 989
rect 162 987 165 989
rect 157 978 165 987
rect 167 989 175 1002
rect 167 987 170 989
rect 172 987 175 989
rect 167 982 175 987
rect 167 980 170 982
rect 172 980 175 982
rect 167 978 175 980
rect 192 989 199 1006
rect 192 987 194 989
rect 196 987 199 989
rect 192 982 199 987
rect 192 980 194 982
rect 196 980 199 982
rect 192 978 199 980
rect 201 978 206 1006
rect 208 978 213 1006
rect 215 996 223 1006
rect 215 994 218 996
rect 220 994 223 996
rect 215 989 223 994
rect 215 987 218 989
rect 220 987 223 989
rect 215 978 223 987
rect 225 978 230 1006
rect 232 978 237 1006
rect 239 989 246 1006
rect 239 987 242 989
rect 244 987 246 989
rect 260 998 267 1000
rect 260 996 262 998
rect 264 996 267 998
rect 260 991 267 996
rect 260 989 262 991
rect 264 989 267 991
rect 260 987 267 989
rect 269 999 274 1000
rect 511 1004 518 1006
rect 293 999 299 1004
rect 269 987 279 999
rect 239 982 246 987
rect 271 986 279 987
rect 281 997 289 999
rect 281 995 284 997
rect 286 995 289 997
rect 281 990 289 995
rect 281 988 284 990
rect 286 988 289 990
rect 281 986 289 988
rect 291 990 299 999
rect 291 988 294 990
rect 296 988 299 990
rect 291 986 299 988
rect 301 1002 308 1004
rect 301 1000 304 1002
rect 306 1000 308 1002
rect 301 995 308 1000
rect 301 993 304 995
rect 306 993 308 995
rect 511 1002 513 1004
rect 515 1002 518 1004
rect 511 997 518 1002
rect 511 995 513 997
rect 515 995 518 997
rect 511 993 518 995
rect 301 991 308 993
rect 301 986 306 991
rect 513 988 518 993
rect 520 989 529 1006
rect 520 988 524 989
rect 239 980 242 982
rect 244 980 246 982
rect 239 978 246 980
rect 271 979 277 986
rect 522 987 524 988
rect 526 987 529 989
rect 522 985 529 987
rect 579 989 586 1005
rect 579 987 581 989
rect 583 987 586 989
rect 579 982 586 987
rect 271 977 273 979
rect 275 977 277 979
rect 271 975 277 977
rect 579 980 581 982
rect 583 980 586 982
rect 579 978 586 980
rect 588 978 593 1005
rect 595 1003 603 1005
rect 595 1001 598 1003
rect 600 1001 603 1003
rect 595 996 603 1001
rect 595 994 598 996
rect 600 994 603 996
rect 595 978 603 994
rect 605 978 610 1005
rect 612 989 619 1005
rect 648 998 654 1005
rect 612 987 615 989
rect 617 987 619 989
rect 612 982 619 987
rect 627 989 634 998
rect 627 987 629 989
rect 631 987 634 989
rect 627 985 634 987
rect 636 996 644 998
rect 636 994 639 996
rect 641 994 644 996
rect 636 989 644 994
rect 636 987 639 989
rect 641 987 644 989
rect 636 985 644 987
rect 646 991 654 998
rect 646 989 649 991
rect 651 989 654 991
rect 646 987 654 989
rect 656 1003 663 1005
rect 656 1001 659 1003
rect 661 1001 663 1003
rect 656 996 663 1001
rect 656 994 659 996
rect 661 994 663 996
rect 656 992 663 994
rect 673 1004 680 1006
rect 673 1002 675 1004
rect 677 1002 680 1004
rect 673 997 680 1002
rect 673 995 675 997
rect 677 995 680 997
rect 673 993 680 995
rect 656 987 661 992
rect 675 988 680 993
rect 682 989 691 1006
rect 682 988 686 989
rect 646 985 652 987
rect 612 980 615 982
rect 617 980 619 982
rect 684 987 686 988
rect 688 987 691 989
rect 684 985 691 987
rect 703 989 710 1005
rect 703 987 705 989
rect 707 987 710 989
rect 703 982 710 987
rect 612 978 619 980
rect 703 980 705 982
rect 707 980 710 982
rect 703 978 710 980
rect 712 978 717 1005
rect 719 1003 727 1005
rect 719 1001 722 1003
rect 724 1001 727 1003
rect 719 996 727 1001
rect 719 994 722 996
rect 724 994 727 996
rect 719 978 727 994
rect 729 978 734 1005
rect 736 989 743 1005
rect 736 987 739 989
rect 741 987 743 989
rect 736 982 743 987
rect 736 980 739 982
rect 741 980 743 982
rect 736 978 743 980
rect 85 959 90 966
rect 83 957 90 959
rect 83 955 85 957
rect 87 955 90 957
rect 83 950 90 955
rect 83 948 85 950
rect 87 948 90 950
rect 83 946 90 948
rect 85 938 90 946
rect 92 938 97 966
rect 99 964 108 966
rect 99 962 104 964
rect 106 962 108 964
rect 99 957 108 962
rect 99 955 104 957
rect 106 955 108 957
rect 127 957 134 959
rect 202 960 207 966
rect 155 957 161 959
rect 127 956 129 957
rect 99 938 108 955
rect 118 951 123 956
rect 116 949 123 951
rect 116 947 118 949
rect 120 947 123 949
rect 116 942 123 947
rect 116 940 118 942
rect 120 940 123 942
rect 116 938 123 940
rect 125 955 129 956
rect 131 955 134 957
rect 125 938 134 955
rect 146 952 151 957
rect 144 950 151 952
rect 144 948 146 950
rect 148 948 151 950
rect 144 943 151 948
rect 144 941 146 943
rect 148 941 151 943
rect 144 939 151 941
rect 153 955 161 957
rect 153 953 156 955
rect 158 953 161 955
rect 153 946 161 953
rect 163 957 171 959
rect 163 955 166 957
rect 168 955 171 957
rect 163 950 171 955
rect 163 948 166 950
rect 168 948 171 950
rect 163 946 171 948
rect 173 957 180 959
rect 173 955 176 957
rect 178 955 180 957
rect 173 946 180 955
rect 200 958 207 960
rect 200 956 202 958
rect 204 956 207 958
rect 200 954 207 956
rect 153 939 159 946
rect 202 939 207 954
rect 209 957 214 966
rect 231 964 243 966
rect 231 962 238 964
rect 240 962 243 964
rect 231 957 243 962
rect 209 950 217 957
rect 209 948 212 950
rect 214 948 217 950
rect 209 939 217 948
rect 219 950 227 957
rect 219 948 222 950
rect 224 948 227 950
rect 219 943 227 948
rect 219 941 222 943
rect 224 941 227 943
rect 219 939 227 941
rect 229 955 238 957
rect 240 955 243 957
rect 229 939 243 955
rect 245 945 250 966
rect 268 957 275 959
rect 268 955 270 957
rect 272 955 275 957
rect 268 946 275 955
rect 277 957 285 959
rect 277 955 280 957
rect 282 955 285 957
rect 277 950 285 955
rect 277 948 280 950
rect 282 948 285 950
rect 277 946 285 948
rect 287 957 293 959
rect 513 960 518 966
rect 511 958 518 960
rect 287 955 295 957
rect 287 953 290 955
rect 292 953 295 955
rect 287 946 295 953
rect 245 943 252 945
rect 245 941 248 943
rect 250 941 252 943
rect 245 939 252 941
rect 289 939 295 946
rect 297 952 302 957
rect 511 956 513 958
rect 515 956 518 958
rect 511 954 518 956
rect 297 950 304 952
rect 297 948 300 950
rect 302 948 304 950
rect 297 943 304 948
rect 297 941 300 943
rect 302 941 304 943
rect 297 939 304 941
rect 513 939 518 954
rect 520 957 525 966
rect 542 964 554 966
rect 542 962 549 964
rect 551 962 554 964
rect 542 957 554 962
rect 520 950 528 957
rect 520 948 523 950
rect 525 948 528 950
rect 520 939 528 948
rect 530 950 538 957
rect 530 948 533 950
rect 535 948 538 950
rect 530 943 538 948
rect 530 941 533 943
rect 535 941 538 943
rect 530 939 538 941
rect 540 955 549 957
rect 551 955 554 957
rect 540 939 554 955
rect 556 945 561 966
rect 590 957 596 959
rect 581 952 586 957
rect 579 950 586 952
rect 579 948 581 950
rect 583 948 586 950
rect 556 943 563 945
rect 579 943 586 948
rect 556 941 559 943
rect 561 941 563 943
rect 556 939 563 941
rect 579 941 581 943
rect 583 941 586 943
rect 579 939 586 941
rect 588 955 596 957
rect 588 953 591 955
rect 593 953 596 955
rect 588 946 596 953
rect 598 957 606 959
rect 598 955 601 957
rect 603 955 606 957
rect 598 950 606 955
rect 598 948 601 950
rect 603 948 606 950
rect 598 946 606 948
rect 608 957 615 959
rect 685 960 690 966
rect 683 958 690 960
rect 608 955 611 957
rect 613 955 615 957
rect 608 946 615 955
rect 623 955 631 957
rect 623 953 626 955
rect 628 953 631 955
rect 588 939 594 946
rect 623 939 631 953
rect 633 950 641 957
rect 633 948 636 950
rect 638 948 641 950
rect 633 943 641 948
rect 633 941 636 943
rect 638 941 641 943
rect 633 939 641 941
rect 643 955 651 957
rect 643 953 646 955
rect 648 953 651 955
rect 643 948 651 953
rect 643 946 646 948
rect 648 946 651 948
rect 643 939 651 946
rect 653 950 661 957
rect 653 948 656 950
rect 658 948 661 950
rect 653 943 661 948
rect 653 941 656 943
rect 658 941 661 943
rect 653 939 661 941
rect 663 955 671 957
rect 663 953 666 955
rect 668 953 671 955
rect 683 956 685 958
rect 687 956 690 958
rect 683 954 690 956
rect 663 948 671 953
rect 663 946 666 948
rect 668 946 671 948
rect 663 939 671 946
rect 685 939 690 954
rect 692 957 697 966
rect 714 964 726 966
rect 714 962 721 964
rect 723 962 726 964
rect 714 957 726 962
rect 692 950 700 957
rect 692 948 695 950
rect 697 948 700 950
rect 692 939 700 948
rect 702 950 710 957
rect 702 948 705 950
rect 707 948 710 950
rect 702 943 710 948
rect 702 941 705 943
rect 707 941 710 943
rect 702 939 710 941
rect 712 955 721 957
rect 723 955 726 957
rect 712 939 726 955
rect 728 945 733 966
rect 728 943 735 945
rect 728 941 731 943
rect 733 941 735 943
rect 728 939 735 941
rect 116 859 123 861
rect 116 857 118 859
rect 120 857 123 859
rect 81 854 89 857
rect 81 852 83 854
rect 85 852 89 854
rect 81 847 89 852
rect 81 845 83 847
rect 85 845 89 847
rect 81 843 89 845
rect 91 854 99 857
rect 91 852 94 854
rect 96 852 99 854
rect 91 847 99 852
rect 91 845 94 847
rect 96 845 99 847
rect 91 843 99 845
rect 101 845 109 857
rect 101 843 105 845
rect 107 843 109 845
rect 116 852 123 857
rect 116 850 118 852
rect 120 850 123 852
rect 116 843 123 850
rect 125 854 131 861
rect 165 859 172 861
rect 165 857 167 859
rect 169 857 172 859
rect 125 847 133 854
rect 125 845 128 847
rect 130 845 133 847
rect 125 843 133 845
rect 103 841 109 843
rect 127 841 133 843
rect 135 852 143 854
rect 135 850 138 852
rect 140 850 143 852
rect 135 845 143 850
rect 135 843 138 845
rect 140 843 143 845
rect 135 841 143 843
rect 145 845 152 854
rect 165 852 172 857
rect 165 850 167 852
rect 169 850 172 852
rect 165 848 172 850
rect 145 843 148 845
rect 150 843 152 845
rect 167 843 172 848
rect 174 854 180 861
rect 239 854 245 861
rect 174 847 182 854
rect 174 845 177 847
rect 179 845 182 847
rect 174 843 182 845
rect 145 841 152 843
rect 176 841 182 843
rect 184 852 192 854
rect 184 850 187 852
rect 189 850 192 852
rect 184 845 192 850
rect 184 843 187 845
rect 189 843 192 845
rect 184 841 192 843
rect 194 845 201 854
rect 194 843 197 845
rect 199 843 201 845
rect 194 841 201 843
rect 218 845 225 854
rect 218 843 220 845
rect 222 843 225 845
rect 218 841 225 843
rect 227 852 235 854
rect 227 850 230 852
rect 232 850 235 852
rect 227 845 235 850
rect 227 843 230 845
rect 232 843 235 845
rect 227 841 235 843
rect 237 847 245 854
rect 237 845 240 847
rect 242 845 245 847
rect 237 843 245 845
rect 247 859 254 861
rect 247 857 250 859
rect 252 857 254 859
rect 247 852 254 857
rect 247 850 250 852
rect 252 850 254 852
rect 247 848 254 850
rect 264 860 271 862
rect 264 858 266 860
rect 268 858 271 860
rect 264 853 271 858
rect 264 851 266 853
rect 268 851 271 853
rect 264 849 271 851
rect 247 843 252 848
rect 266 844 271 849
rect 273 845 282 862
rect 292 859 299 861
rect 292 857 294 859
rect 296 857 299 859
rect 292 852 299 857
rect 292 850 294 852
rect 296 850 299 852
rect 292 848 299 850
rect 273 844 277 845
rect 237 841 243 843
rect 275 843 277 844
rect 279 843 282 845
rect 294 843 299 848
rect 301 854 307 861
rect 336 858 343 860
rect 336 856 338 858
rect 340 856 343 858
rect 301 847 309 854
rect 301 845 304 847
rect 306 845 309 847
rect 301 843 309 845
rect 275 841 282 843
rect 303 841 309 843
rect 311 852 319 854
rect 311 850 314 852
rect 316 850 319 852
rect 311 845 319 850
rect 311 843 314 845
rect 316 843 319 845
rect 311 841 319 843
rect 321 845 328 854
rect 336 851 343 856
rect 336 849 338 851
rect 340 849 343 851
rect 336 847 343 849
rect 321 843 324 845
rect 326 843 328 845
rect 321 841 328 843
rect 338 842 343 847
rect 345 855 351 860
rect 370 855 375 856
rect 345 846 353 855
rect 345 844 348 846
rect 350 844 353 846
rect 345 842 353 844
rect 355 853 363 855
rect 355 851 358 853
rect 360 851 363 853
rect 355 846 363 851
rect 355 844 358 846
rect 360 844 363 846
rect 355 842 363 844
rect 365 843 375 855
rect 377 854 384 856
rect 507 854 513 861
rect 377 852 380 854
rect 382 852 384 854
rect 377 847 384 852
rect 377 845 380 847
rect 382 845 384 847
rect 377 843 384 845
rect 486 845 493 854
rect 486 843 488 845
rect 490 843 493 845
rect 365 842 373 843
rect 367 835 373 842
rect 486 841 493 843
rect 495 852 503 854
rect 495 850 498 852
rect 500 850 503 852
rect 495 845 503 850
rect 495 843 498 845
rect 500 843 503 845
rect 495 841 503 843
rect 505 847 513 854
rect 505 845 508 847
rect 510 845 513 847
rect 505 843 513 845
rect 515 859 522 861
rect 515 857 518 859
rect 520 857 522 859
rect 515 852 522 857
rect 515 850 518 852
rect 520 850 522 852
rect 515 848 522 850
rect 531 860 538 862
rect 531 858 533 860
rect 535 858 538 860
rect 531 853 538 858
rect 531 851 533 853
rect 535 851 538 853
rect 531 849 538 851
rect 515 843 520 848
rect 533 844 538 849
rect 540 845 549 862
rect 580 854 586 861
rect 540 844 544 845
rect 505 841 511 843
rect 367 833 369 835
rect 371 833 373 835
rect 367 831 373 833
rect 542 843 544 844
rect 546 843 549 845
rect 542 841 549 843
rect 559 845 566 854
rect 559 843 561 845
rect 563 843 566 845
rect 559 841 566 843
rect 568 852 576 854
rect 568 850 571 852
rect 573 850 576 852
rect 568 845 576 850
rect 568 843 571 845
rect 573 843 576 845
rect 568 841 576 843
rect 578 847 586 854
rect 578 845 581 847
rect 583 845 586 847
rect 578 843 586 845
rect 588 859 595 861
rect 588 857 591 859
rect 593 857 595 859
rect 588 852 595 857
rect 588 850 591 852
rect 593 850 595 852
rect 588 848 595 850
rect 607 859 614 861
rect 607 857 609 859
rect 611 857 614 859
rect 607 852 614 857
rect 607 850 609 852
rect 611 850 614 852
rect 607 848 614 850
rect 588 843 593 848
rect 609 843 614 848
rect 616 854 622 861
rect 651 854 658 856
rect 616 847 624 854
rect 616 845 619 847
rect 621 845 624 847
rect 616 843 624 845
rect 578 841 584 843
rect 618 841 624 843
rect 626 852 634 854
rect 626 850 629 852
rect 631 850 634 852
rect 626 845 634 850
rect 626 843 629 845
rect 631 843 634 845
rect 626 841 634 843
rect 636 845 643 854
rect 636 843 639 845
rect 641 843 643 845
rect 651 852 653 854
rect 655 852 658 854
rect 651 847 658 852
rect 651 845 653 847
rect 655 845 658 847
rect 651 843 658 845
rect 660 855 665 856
rect 684 855 690 860
rect 660 843 670 855
rect 636 841 643 843
rect 662 842 670 843
rect 672 853 680 855
rect 672 851 675 853
rect 677 851 680 853
rect 672 846 680 851
rect 672 844 675 846
rect 677 844 680 846
rect 672 842 680 844
rect 682 846 690 855
rect 682 844 685 846
rect 687 844 690 846
rect 682 842 690 844
rect 692 858 699 860
rect 692 856 695 858
rect 697 856 699 858
rect 692 851 699 856
rect 692 849 695 851
rect 697 849 699 851
rect 692 847 699 849
rect 692 842 697 847
rect 707 845 714 854
rect 707 843 709 845
rect 711 843 714 845
rect 662 835 668 842
rect 707 838 714 843
rect 662 833 664 835
rect 666 833 668 835
rect 707 836 709 838
rect 711 836 714 838
rect 707 834 714 836
rect 716 852 724 854
rect 716 850 719 852
rect 721 850 724 852
rect 716 845 724 850
rect 716 843 719 845
rect 721 843 724 845
rect 716 834 724 843
rect 726 845 734 854
rect 726 843 729 845
rect 731 843 734 845
rect 726 838 734 843
rect 726 836 729 838
rect 731 836 734 838
rect 726 834 734 836
rect 736 852 743 854
rect 736 850 739 852
rect 741 850 743 852
rect 736 845 743 850
rect 736 843 739 845
rect 741 843 743 845
rect 736 841 743 843
rect 736 834 741 841
rect 662 831 668 833
rect 155 823 161 825
rect 82 815 87 822
rect 80 813 87 815
rect 80 811 82 813
rect 84 811 87 813
rect 80 806 87 811
rect 80 804 82 806
rect 84 804 87 806
rect 80 802 87 804
rect 89 820 97 822
rect 89 818 92 820
rect 94 818 97 820
rect 89 813 97 818
rect 89 811 92 813
rect 94 811 97 813
rect 89 802 97 811
rect 99 813 107 822
rect 99 811 102 813
rect 104 811 107 813
rect 99 806 107 811
rect 99 804 102 806
rect 104 804 107 806
rect 99 802 107 804
rect 109 820 116 822
rect 109 818 112 820
rect 114 818 116 820
rect 155 821 157 823
rect 159 821 161 823
rect 109 813 116 818
rect 155 814 161 821
rect 109 811 112 813
rect 114 811 116 813
rect 109 802 116 811
rect 126 809 131 814
rect 124 807 131 809
rect 124 805 126 807
rect 128 805 131 807
rect 124 800 131 805
rect 124 798 126 800
rect 128 798 131 800
rect 124 796 131 798
rect 133 812 141 814
rect 133 810 136 812
rect 138 810 141 812
rect 133 801 141 810
rect 143 812 151 814
rect 143 810 146 812
rect 148 810 151 812
rect 143 805 151 810
rect 143 803 146 805
rect 148 803 151 805
rect 143 801 151 803
rect 153 813 161 814
rect 180 813 187 815
rect 153 801 163 813
rect 133 796 139 801
rect 158 800 163 801
rect 165 811 172 813
rect 165 809 168 811
rect 170 809 172 811
rect 165 804 172 809
rect 165 802 168 804
rect 170 802 172 804
rect 180 811 182 813
rect 184 811 187 813
rect 180 802 187 811
rect 189 813 197 815
rect 189 811 192 813
rect 194 811 197 813
rect 189 806 197 811
rect 189 804 192 806
rect 194 804 197 806
rect 189 802 197 804
rect 199 813 205 815
rect 239 813 245 815
rect 199 811 207 813
rect 199 809 202 811
rect 204 809 207 811
rect 199 802 207 809
rect 165 800 172 802
rect 201 795 207 802
rect 209 808 214 813
rect 230 808 235 813
rect 209 806 216 808
rect 209 804 212 806
rect 214 804 216 806
rect 209 799 216 804
rect 209 797 212 799
rect 214 797 216 799
rect 209 795 216 797
rect 228 806 235 808
rect 228 804 230 806
rect 232 804 235 806
rect 228 799 235 804
rect 228 797 230 799
rect 232 797 235 799
rect 228 795 235 797
rect 237 811 245 813
rect 237 809 240 811
rect 242 809 245 811
rect 237 802 245 809
rect 247 813 255 815
rect 247 811 250 813
rect 252 811 255 813
rect 247 806 255 811
rect 247 804 250 806
rect 252 804 255 806
rect 247 802 255 804
rect 257 813 264 815
rect 257 811 260 813
rect 262 811 264 813
rect 257 802 264 811
rect 274 813 281 815
rect 274 811 277 813
rect 279 812 281 813
rect 450 823 456 825
rect 450 821 452 823
rect 454 821 456 823
rect 312 813 318 815
rect 279 811 283 812
rect 237 795 243 802
rect 274 794 283 811
rect 285 807 290 812
rect 303 808 308 813
rect 285 805 292 807
rect 285 803 288 805
rect 290 803 292 805
rect 285 798 292 803
rect 285 796 288 798
rect 290 796 292 798
rect 285 794 292 796
rect 301 806 308 808
rect 301 804 303 806
rect 305 804 308 806
rect 301 799 308 804
rect 301 797 303 799
rect 305 797 308 799
rect 301 795 308 797
rect 310 811 318 813
rect 310 809 313 811
rect 315 809 318 811
rect 310 802 318 809
rect 320 813 328 815
rect 320 811 323 813
rect 325 811 328 813
rect 320 806 328 811
rect 320 804 323 806
rect 325 804 328 806
rect 320 802 328 804
rect 330 813 337 815
rect 450 814 456 821
rect 450 813 458 814
rect 330 811 333 813
rect 335 811 337 813
rect 330 802 337 811
rect 439 811 446 813
rect 439 809 441 811
rect 443 809 446 811
rect 439 804 446 809
rect 439 802 441 804
rect 443 802 446 804
rect 310 795 316 802
rect 439 800 446 802
rect 448 801 458 813
rect 460 812 468 814
rect 460 810 463 812
rect 465 810 468 812
rect 460 805 468 810
rect 460 803 463 805
rect 465 803 468 805
rect 460 801 468 803
rect 470 812 478 814
rect 470 810 473 812
rect 475 810 478 812
rect 470 801 478 810
rect 448 800 453 801
rect 472 796 478 801
rect 480 809 485 814
rect 495 813 502 815
rect 495 811 497 813
rect 499 811 502 813
rect 480 807 487 809
rect 480 805 483 807
rect 485 805 487 807
rect 480 800 487 805
rect 495 802 502 811
rect 504 813 512 815
rect 504 811 507 813
rect 509 811 512 813
rect 504 806 512 811
rect 504 804 507 806
rect 509 804 512 806
rect 504 802 512 804
rect 514 813 520 815
rect 541 813 548 815
rect 514 811 522 813
rect 514 809 517 811
rect 519 809 522 811
rect 514 802 522 809
rect 480 798 483 800
rect 485 798 487 800
rect 480 796 487 798
rect 516 795 522 802
rect 524 808 529 813
rect 541 811 544 813
rect 546 812 548 813
rect 580 813 586 815
rect 546 811 550 812
rect 524 806 531 808
rect 524 804 527 806
rect 529 804 531 806
rect 524 799 531 804
rect 524 797 527 799
rect 529 797 531 799
rect 524 795 531 797
rect 541 794 550 811
rect 552 807 557 812
rect 571 808 576 813
rect 552 805 559 807
rect 552 803 555 805
rect 557 803 559 805
rect 552 798 559 803
rect 552 796 555 798
rect 557 796 559 798
rect 552 794 559 796
rect 569 806 576 808
rect 569 804 571 806
rect 573 804 576 806
rect 569 799 576 804
rect 569 797 571 799
rect 573 797 576 799
rect 569 795 576 797
rect 578 811 586 813
rect 578 809 581 811
rect 583 809 586 811
rect 578 802 586 809
rect 588 813 596 815
rect 588 811 591 813
rect 593 811 596 813
rect 588 806 596 811
rect 588 804 591 806
rect 593 804 596 806
rect 588 802 596 804
rect 598 813 605 815
rect 598 811 601 813
rect 603 811 605 813
rect 598 802 605 811
rect 622 813 629 815
rect 622 811 624 813
rect 626 811 629 813
rect 622 802 629 811
rect 631 813 639 815
rect 631 811 634 813
rect 636 811 639 813
rect 631 806 639 811
rect 631 804 634 806
rect 636 804 639 806
rect 631 802 639 804
rect 641 813 647 815
rect 671 813 678 815
rect 641 811 649 813
rect 641 809 644 811
rect 646 809 649 811
rect 641 802 649 809
rect 578 795 584 802
rect 643 795 649 802
rect 651 808 656 813
rect 671 811 673 813
rect 675 811 678 813
rect 651 806 658 808
rect 651 804 654 806
rect 656 804 658 806
rect 651 799 658 804
rect 671 802 678 811
rect 680 813 688 815
rect 680 811 683 813
rect 685 811 688 813
rect 680 806 688 811
rect 680 804 683 806
rect 685 804 688 806
rect 680 802 688 804
rect 690 813 696 815
rect 714 813 720 815
rect 690 811 698 813
rect 690 809 693 811
rect 695 809 698 811
rect 690 802 698 809
rect 651 797 654 799
rect 656 797 658 799
rect 651 795 658 797
rect 692 795 698 802
rect 700 806 707 813
rect 700 804 703 806
rect 705 804 707 806
rect 700 799 707 804
rect 714 811 716 813
rect 718 811 722 813
rect 714 799 722 811
rect 724 811 732 813
rect 724 809 727 811
rect 729 809 732 811
rect 724 804 732 809
rect 724 802 727 804
rect 729 802 732 804
rect 724 799 732 802
rect 734 811 742 813
rect 734 809 738 811
rect 740 809 742 811
rect 734 804 742 809
rect 734 802 738 804
rect 740 802 742 804
rect 734 799 742 802
rect 700 797 703 799
rect 705 797 707 799
rect 700 795 707 797
rect 88 715 95 717
rect 88 713 90 715
rect 92 713 95 715
rect 88 711 95 713
rect 90 690 95 711
rect 97 701 111 717
rect 97 699 100 701
rect 102 699 111 701
rect 113 715 121 717
rect 113 713 116 715
rect 118 713 121 715
rect 113 708 121 713
rect 113 706 116 708
rect 118 706 121 708
rect 113 699 121 706
rect 123 708 131 717
rect 123 706 126 708
rect 128 706 131 708
rect 123 699 131 706
rect 97 694 109 699
rect 97 692 100 694
rect 102 692 109 694
rect 97 690 109 692
rect 126 690 131 699
rect 133 702 138 717
rect 152 710 160 717
rect 152 708 155 710
rect 157 708 160 710
rect 152 703 160 708
rect 133 700 140 702
rect 133 698 136 700
rect 138 698 140 700
rect 152 701 155 703
rect 157 701 160 703
rect 152 699 160 701
rect 162 715 170 717
rect 162 713 165 715
rect 167 713 170 715
rect 162 708 170 713
rect 162 706 165 708
rect 167 706 170 708
rect 162 699 170 706
rect 172 710 180 717
rect 172 708 175 710
rect 177 708 180 710
rect 172 703 180 708
rect 172 701 175 703
rect 177 701 180 703
rect 172 699 180 701
rect 182 715 190 717
rect 182 713 185 715
rect 187 713 190 715
rect 182 708 190 713
rect 182 706 185 708
rect 187 706 190 708
rect 182 699 190 706
rect 192 703 200 717
rect 229 710 235 717
rect 192 701 195 703
rect 197 701 200 703
rect 192 699 200 701
rect 208 701 215 710
rect 208 699 210 701
rect 212 699 215 701
rect 133 696 140 698
rect 133 690 138 696
rect 208 697 215 699
rect 217 708 225 710
rect 217 706 220 708
rect 222 706 225 708
rect 217 701 225 706
rect 217 699 220 701
rect 222 699 225 701
rect 217 697 225 699
rect 227 703 235 710
rect 227 701 230 703
rect 232 701 235 703
rect 227 699 235 701
rect 237 715 244 717
rect 237 713 240 715
rect 242 713 244 715
rect 260 715 267 717
rect 260 713 262 715
rect 264 713 267 715
rect 237 708 244 713
rect 260 711 267 713
rect 237 706 240 708
rect 242 706 244 708
rect 237 704 244 706
rect 237 699 242 704
rect 227 697 233 699
rect 262 690 267 711
rect 269 701 283 717
rect 269 699 272 701
rect 274 699 283 701
rect 285 715 293 717
rect 285 713 288 715
rect 290 713 293 715
rect 285 708 293 713
rect 285 706 288 708
rect 290 706 293 708
rect 285 699 293 706
rect 295 708 303 717
rect 295 706 298 708
rect 300 706 303 708
rect 295 699 303 706
rect 269 694 281 699
rect 269 692 272 694
rect 274 692 281 694
rect 269 690 281 692
rect 298 690 303 699
rect 305 702 310 717
rect 320 716 327 718
rect 320 714 322 716
rect 324 714 327 716
rect 320 709 327 714
rect 320 707 322 709
rect 324 707 327 709
rect 320 705 327 707
rect 305 700 312 702
rect 322 700 327 705
rect 329 701 338 718
rect 519 715 526 717
rect 519 713 521 715
rect 523 713 526 715
rect 519 708 526 713
rect 519 706 521 708
rect 523 706 526 708
rect 519 704 526 706
rect 329 700 333 701
rect 305 698 308 700
rect 310 698 312 700
rect 305 696 312 698
rect 305 690 310 696
rect 331 699 333 700
rect 335 699 338 701
rect 521 699 526 704
rect 528 710 534 717
rect 571 715 578 717
rect 571 713 573 715
rect 575 713 578 715
rect 571 711 578 713
rect 528 703 536 710
rect 528 701 531 703
rect 533 701 536 703
rect 528 699 536 701
rect 331 697 338 699
rect 530 697 536 699
rect 538 708 546 710
rect 538 706 541 708
rect 543 706 546 708
rect 538 701 546 706
rect 538 699 541 701
rect 543 699 546 701
rect 538 697 546 699
rect 548 701 555 710
rect 548 699 551 701
rect 553 699 555 701
rect 548 697 555 699
rect 573 690 578 711
rect 580 701 594 717
rect 580 699 583 701
rect 585 699 594 701
rect 596 715 604 717
rect 596 713 599 715
rect 601 713 604 715
rect 596 708 604 713
rect 596 706 599 708
rect 601 706 604 708
rect 596 699 604 706
rect 606 708 614 717
rect 606 706 609 708
rect 611 706 614 708
rect 606 699 614 706
rect 580 694 592 699
rect 580 692 583 694
rect 585 692 592 694
rect 580 690 592 692
rect 609 690 614 699
rect 616 702 621 717
rect 664 710 670 717
rect 616 700 623 702
rect 616 698 619 700
rect 621 698 623 700
rect 616 696 623 698
rect 643 701 650 710
rect 643 699 645 701
rect 647 699 650 701
rect 643 697 650 699
rect 652 708 660 710
rect 652 706 655 708
rect 657 706 660 708
rect 652 701 660 706
rect 652 699 655 701
rect 657 699 660 701
rect 652 697 660 699
rect 662 703 670 710
rect 662 701 665 703
rect 667 701 670 703
rect 662 699 670 701
rect 672 715 679 717
rect 672 713 675 715
rect 677 713 679 715
rect 672 708 679 713
rect 672 706 675 708
rect 677 706 679 708
rect 672 704 679 706
rect 672 699 677 704
rect 689 701 698 718
rect 689 699 692 701
rect 694 700 698 701
rect 700 716 707 718
rect 700 714 703 716
rect 705 714 707 716
rect 700 709 707 714
rect 700 707 703 709
rect 705 707 707 709
rect 700 705 707 707
rect 700 700 705 705
rect 715 701 724 718
rect 694 699 696 700
rect 662 697 668 699
rect 616 690 621 696
rect 689 697 696 699
rect 715 699 717 701
rect 719 699 724 701
rect 715 694 724 699
rect 715 692 717 694
rect 719 692 724 694
rect 715 690 724 692
rect 726 690 731 718
rect 733 710 738 718
rect 733 708 740 710
rect 733 706 736 708
rect 738 706 740 708
rect 733 701 740 706
rect 733 699 736 701
rect 738 699 740 701
rect 733 697 740 699
rect 733 690 738 697
rect 80 676 87 678
rect 80 674 82 676
rect 84 674 87 676
rect 80 669 87 674
rect 80 667 82 669
rect 84 667 87 669
rect 80 651 87 667
rect 89 651 94 678
rect 96 662 104 678
rect 96 660 99 662
rect 101 660 104 662
rect 96 655 104 660
rect 96 653 99 655
rect 101 653 104 655
rect 96 651 104 653
rect 106 651 111 678
rect 113 676 120 678
rect 113 674 116 676
rect 118 674 120 676
rect 546 679 552 681
rect 204 676 211 678
rect 113 669 120 674
rect 113 667 116 669
rect 118 667 120 669
rect 113 651 120 667
rect 132 669 139 671
rect 132 667 135 669
rect 137 668 139 669
rect 204 674 206 676
rect 208 674 211 676
rect 171 669 177 671
rect 137 667 141 668
rect 132 650 141 667
rect 143 663 148 668
rect 162 664 167 669
rect 143 661 150 663
rect 143 659 146 661
rect 148 659 150 661
rect 143 654 150 659
rect 143 652 146 654
rect 148 652 150 654
rect 143 650 150 652
rect 160 662 167 664
rect 160 660 162 662
rect 164 660 167 662
rect 160 655 167 660
rect 160 653 162 655
rect 164 653 167 655
rect 160 651 167 653
rect 169 667 177 669
rect 169 665 172 667
rect 174 665 177 667
rect 169 658 177 665
rect 179 669 187 671
rect 179 667 182 669
rect 184 667 187 669
rect 179 662 187 667
rect 179 660 182 662
rect 184 660 187 662
rect 179 658 187 660
rect 189 669 196 671
rect 189 667 192 669
rect 194 667 196 669
rect 189 658 196 667
rect 204 669 211 674
rect 204 667 206 669
rect 208 667 211 669
rect 169 651 175 658
rect 204 651 211 667
rect 213 651 218 678
rect 220 662 228 678
rect 220 660 223 662
rect 225 660 228 662
rect 220 655 228 660
rect 220 653 223 655
rect 225 653 228 655
rect 220 651 228 653
rect 230 651 235 678
rect 237 676 244 678
rect 237 674 240 676
rect 242 674 244 676
rect 546 677 548 679
rect 550 677 552 679
rect 237 669 244 674
rect 546 670 552 677
rect 577 676 584 678
rect 577 674 579 676
rect 581 674 584 676
rect 237 667 240 669
rect 242 667 244 669
rect 237 651 244 667
rect 517 665 522 670
rect 515 663 522 665
rect 515 661 517 663
rect 519 661 522 663
rect 515 656 522 661
rect 515 654 517 656
rect 519 654 522 656
rect 515 652 522 654
rect 524 668 532 670
rect 524 666 527 668
rect 529 666 532 668
rect 524 657 532 666
rect 534 668 542 670
rect 534 666 537 668
rect 539 666 542 668
rect 534 661 542 666
rect 534 659 537 661
rect 539 659 542 661
rect 534 657 542 659
rect 544 669 552 670
rect 577 669 584 674
rect 544 657 554 669
rect 524 652 530 657
rect 549 656 554 657
rect 556 667 563 669
rect 556 665 559 667
rect 561 665 563 667
rect 556 660 563 665
rect 556 658 559 660
rect 561 658 563 660
rect 556 656 563 658
rect 577 667 579 669
rect 581 667 584 669
rect 577 650 584 667
rect 586 650 591 678
rect 593 650 598 678
rect 600 669 608 678
rect 600 667 603 669
rect 605 667 608 669
rect 600 662 608 667
rect 600 660 603 662
rect 605 660 608 662
rect 600 650 608 660
rect 610 650 615 678
rect 617 650 622 678
rect 624 676 631 678
rect 624 674 627 676
rect 629 674 631 676
rect 624 669 631 674
rect 624 667 627 669
rect 629 667 631 669
rect 624 650 631 667
rect 648 676 656 678
rect 648 674 651 676
rect 653 674 656 676
rect 648 669 656 674
rect 648 667 651 669
rect 653 667 656 669
rect 648 654 656 667
rect 658 669 666 678
rect 658 667 661 669
rect 663 667 666 669
rect 658 662 666 667
rect 658 660 661 662
rect 663 660 666 662
rect 658 654 666 660
rect 668 676 675 678
rect 668 674 671 676
rect 673 674 675 676
rect 668 669 675 674
rect 685 672 690 678
rect 668 667 671 669
rect 673 667 675 669
rect 668 654 675 667
rect 683 670 690 672
rect 683 668 685 670
rect 687 668 690 670
rect 683 666 690 668
rect 685 651 690 666
rect 692 669 697 678
rect 714 676 726 678
rect 714 674 721 676
rect 723 674 726 676
rect 714 669 726 674
rect 692 662 700 669
rect 692 660 695 662
rect 697 660 700 662
rect 692 651 700 660
rect 702 662 710 669
rect 702 660 705 662
rect 707 660 710 662
rect 702 655 710 660
rect 702 653 705 655
rect 707 653 710 655
rect 702 651 710 653
rect 712 667 721 669
rect 723 667 726 669
rect 712 651 726 667
rect 728 657 733 678
rect 728 655 735 657
rect 728 653 731 655
rect 733 653 735 655
rect 728 651 735 653
rect 88 571 95 573
rect 88 569 90 571
rect 92 569 95 571
rect 88 567 95 569
rect 90 546 95 567
rect 97 557 111 573
rect 97 555 100 557
rect 102 555 111 557
rect 113 571 121 573
rect 113 569 116 571
rect 118 569 121 571
rect 113 564 121 569
rect 113 562 116 564
rect 118 562 121 564
rect 113 555 121 562
rect 123 564 131 573
rect 123 562 126 564
rect 128 562 131 564
rect 123 555 131 562
rect 97 550 109 555
rect 97 548 100 550
rect 102 548 109 550
rect 97 546 109 548
rect 126 546 131 555
rect 133 558 138 573
rect 133 556 140 558
rect 133 554 136 556
rect 138 554 140 556
rect 133 552 140 554
rect 148 557 155 570
rect 148 555 150 557
rect 152 555 155 557
rect 133 546 138 552
rect 148 550 155 555
rect 148 548 150 550
rect 152 548 155 550
rect 148 546 155 548
rect 157 564 165 570
rect 157 562 160 564
rect 162 562 165 564
rect 157 557 165 562
rect 157 555 160 557
rect 162 555 165 557
rect 157 546 165 555
rect 167 557 175 570
rect 207 566 213 573
rect 167 555 170 557
rect 172 555 175 557
rect 167 550 175 555
rect 186 557 193 566
rect 186 555 188 557
rect 190 555 193 557
rect 186 553 193 555
rect 195 564 203 566
rect 195 562 198 564
rect 200 562 203 564
rect 195 557 203 562
rect 195 555 198 557
rect 200 555 203 557
rect 195 553 203 555
rect 205 559 213 566
rect 205 557 208 559
rect 210 557 213 559
rect 205 555 213 557
rect 215 571 222 573
rect 215 569 218 571
rect 220 569 222 571
rect 215 564 222 569
rect 215 562 218 564
rect 220 562 222 564
rect 215 560 222 562
rect 234 572 241 574
rect 234 570 236 572
rect 238 570 241 572
rect 234 565 241 570
rect 234 563 236 565
rect 238 563 241 565
rect 234 561 241 563
rect 215 555 220 560
rect 236 556 241 561
rect 243 557 252 574
rect 243 556 247 557
rect 205 553 211 555
rect 167 548 170 550
rect 172 548 175 550
rect 245 555 247 556
rect 249 555 252 557
rect 495 566 502 573
rect 495 564 497 566
rect 499 564 502 566
rect 495 559 502 564
rect 495 557 497 559
rect 499 557 502 559
rect 495 555 502 557
rect 504 555 509 573
rect 511 555 516 573
rect 518 555 523 573
rect 525 565 533 573
rect 525 563 528 565
rect 530 563 533 565
rect 525 555 533 563
rect 245 553 252 555
rect 167 546 175 548
rect 528 548 533 555
rect 535 548 540 573
rect 542 548 547 573
rect 549 548 554 573
rect 556 548 565 573
rect 587 566 594 568
rect 587 564 589 566
rect 591 564 594 566
rect 587 559 594 564
rect 587 557 589 559
rect 591 557 594 559
rect 587 555 594 557
rect 596 567 601 568
rect 620 567 626 572
rect 596 555 606 567
rect 598 554 606 555
rect 608 565 616 567
rect 608 563 611 565
rect 613 563 616 565
rect 608 558 616 563
rect 608 556 611 558
rect 613 556 616 558
rect 608 554 616 556
rect 618 558 626 567
rect 618 556 621 558
rect 623 556 626 558
rect 618 554 626 556
rect 628 570 635 572
rect 628 568 631 570
rect 633 568 635 570
rect 628 563 635 568
rect 664 566 670 573
rect 628 561 631 563
rect 633 561 635 563
rect 628 559 635 561
rect 628 554 633 559
rect 643 557 650 566
rect 643 555 645 557
rect 647 555 650 557
rect 558 547 565 548
rect 558 545 560 547
rect 562 545 565 547
rect 558 543 565 545
rect 598 547 604 554
rect 643 553 650 555
rect 652 564 660 566
rect 652 562 655 564
rect 657 562 660 564
rect 652 557 660 562
rect 652 555 655 557
rect 657 555 660 557
rect 652 553 660 555
rect 662 559 670 566
rect 662 557 665 559
rect 667 557 670 559
rect 662 555 670 557
rect 672 571 679 573
rect 672 569 675 571
rect 677 569 679 571
rect 672 564 679 569
rect 672 562 675 564
rect 677 562 679 564
rect 672 560 679 562
rect 672 555 677 560
rect 689 557 698 574
rect 689 555 692 557
rect 694 556 698 557
rect 700 572 707 574
rect 700 570 703 572
rect 705 570 707 572
rect 700 565 707 570
rect 700 563 703 565
rect 705 563 707 565
rect 700 561 707 563
rect 700 556 705 561
rect 716 557 724 570
rect 694 555 696 556
rect 662 553 668 555
rect 689 553 696 555
rect 716 555 719 557
rect 721 555 724 557
rect 716 550 724 555
rect 598 545 600 547
rect 602 545 604 547
rect 598 543 604 545
rect 716 548 719 550
rect 721 548 724 550
rect 716 546 724 548
rect 726 564 734 570
rect 726 562 729 564
rect 731 562 734 564
rect 726 557 734 562
rect 726 555 729 557
rect 731 555 734 557
rect 726 546 734 555
rect 736 557 743 570
rect 736 555 739 557
rect 741 555 743 557
rect 736 550 743 555
rect 736 548 739 550
rect 741 548 743 550
rect 736 546 743 548
rect 80 532 87 534
rect 80 530 82 532
rect 84 530 87 532
rect 80 525 87 530
rect 80 523 82 525
rect 84 523 87 525
rect 80 507 87 523
rect 89 507 94 534
rect 96 518 104 534
rect 96 516 99 518
rect 101 516 104 518
rect 96 511 104 516
rect 96 509 99 511
rect 101 509 104 511
rect 96 507 104 509
rect 106 507 111 534
rect 113 532 120 534
rect 113 530 116 532
rect 118 530 120 532
rect 113 525 120 530
rect 113 523 116 525
rect 118 523 120 525
rect 113 507 120 523
rect 130 525 137 527
rect 130 523 133 525
rect 135 524 137 525
rect 161 528 166 534
rect 159 526 166 528
rect 159 524 161 526
rect 163 524 166 526
rect 135 523 139 524
rect 130 506 139 523
rect 141 519 146 524
rect 159 522 166 524
rect 141 517 148 519
rect 141 515 144 517
rect 146 515 148 517
rect 141 510 148 515
rect 141 508 144 510
rect 146 508 148 510
rect 141 506 148 508
rect 161 507 166 522
rect 168 525 173 534
rect 190 532 202 534
rect 190 530 197 532
rect 199 530 202 532
rect 190 525 202 530
rect 168 518 176 525
rect 168 516 171 518
rect 173 516 176 518
rect 168 507 176 516
rect 178 518 186 525
rect 178 516 181 518
rect 183 516 186 518
rect 178 511 186 516
rect 178 509 181 511
rect 183 509 186 511
rect 178 507 186 509
rect 188 523 197 525
rect 199 523 202 525
rect 188 507 202 523
rect 204 513 209 534
rect 242 525 247 533
rect 229 523 237 525
rect 229 521 232 523
rect 234 521 237 523
rect 229 516 237 521
rect 229 514 232 516
rect 234 514 237 516
rect 204 511 211 513
rect 204 509 207 511
rect 209 509 211 511
rect 204 507 211 509
rect 229 509 237 514
rect 239 517 247 525
rect 239 515 242 517
rect 244 515 247 517
rect 239 509 247 515
rect 249 531 257 533
rect 478 535 484 537
rect 478 533 480 535
rect 482 533 484 535
rect 249 529 252 531
rect 254 529 257 531
rect 478 530 484 533
rect 249 524 257 529
rect 249 522 252 524
rect 254 522 257 524
rect 249 509 257 522
rect 447 525 454 527
rect 447 523 450 525
rect 452 524 454 525
rect 452 523 456 524
rect 447 506 456 523
rect 458 519 463 524
rect 458 517 465 519
rect 458 515 461 517
rect 463 515 465 517
rect 458 510 465 515
rect 478 513 486 530
rect 488 525 496 530
rect 488 523 491 525
rect 493 523 496 525
rect 488 518 496 523
rect 488 516 491 518
rect 493 516 496 518
rect 488 513 496 516
rect 498 528 506 530
rect 498 526 501 528
rect 503 526 506 528
rect 498 513 506 526
rect 508 525 516 530
rect 508 523 511 525
rect 513 523 516 525
rect 508 518 516 523
rect 508 516 511 518
rect 513 516 516 518
rect 508 513 516 516
rect 518 528 525 530
rect 537 528 542 534
rect 518 526 521 528
rect 523 526 525 528
rect 518 513 525 526
rect 535 526 542 528
rect 535 524 537 526
rect 539 524 542 526
rect 535 522 542 524
rect 458 508 461 510
rect 463 508 465 510
rect 458 506 465 508
rect 537 507 542 522
rect 544 525 549 534
rect 566 532 578 534
rect 566 530 573 532
rect 575 530 578 532
rect 566 525 578 530
rect 544 518 552 525
rect 544 516 547 518
rect 549 516 552 518
rect 544 507 552 516
rect 554 518 562 525
rect 554 516 557 518
rect 559 516 562 518
rect 554 511 562 516
rect 554 509 557 511
rect 559 509 562 511
rect 554 507 562 509
rect 564 523 573 525
rect 575 523 578 525
rect 564 507 578 523
rect 580 513 585 534
rect 647 532 656 534
rect 647 530 649 532
rect 651 530 656 532
rect 603 525 610 527
rect 603 523 605 525
rect 607 523 610 525
rect 603 514 610 523
rect 612 525 620 527
rect 612 523 615 525
rect 617 523 620 525
rect 612 518 620 523
rect 612 516 615 518
rect 617 516 620 518
rect 612 514 620 516
rect 622 525 628 527
rect 647 525 656 530
rect 622 523 630 525
rect 622 521 625 523
rect 627 521 630 523
rect 622 514 630 521
rect 580 511 587 513
rect 580 509 583 511
rect 585 509 587 511
rect 580 507 587 509
rect 624 507 630 514
rect 632 520 637 525
rect 647 523 649 525
rect 651 523 656 525
rect 632 518 639 520
rect 632 516 635 518
rect 637 516 639 518
rect 632 511 639 516
rect 632 509 635 511
rect 637 509 639 511
rect 632 507 639 509
rect 647 506 656 523
rect 658 506 663 534
rect 665 527 670 534
rect 685 528 690 534
rect 665 525 672 527
rect 665 523 668 525
rect 670 523 672 525
rect 665 518 672 523
rect 683 526 690 528
rect 683 524 685 526
rect 687 524 690 526
rect 683 522 690 524
rect 665 516 668 518
rect 670 516 672 518
rect 665 514 672 516
rect 665 506 670 514
rect 685 507 690 522
rect 692 525 697 534
rect 714 532 726 534
rect 714 530 721 532
rect 723 530 726 532
rect 714 525 726 530
rect 692 518 700 525
rect 692 516 695 518
rect 697 516 700 518
rect 692 507 700 516
rect 702 518 710 525
rect 702 516 705 518
rect 707 516 710 518
rect 702 511 710 516
rect 702 509 705 511
rect 707 509 710 511
rect 702 507 710 509
rect 712 523 721 525
rect 723 523 726 525
rect 712 507 726 523
rect 728 513 733 534
rect 728 511 735 513
rect 728 509 731 511
rect 733 509 735 511
rect 728 507 735 509
rect 7 320 12 327
rect 5 318 12 320
rect 5 316 7 318
rect 9 316 12 318
rect 5 314 12 316
rect 14 314 23 327
rect 16 310 23 314
rect 16 308 18 310
rect 20 308 23 310
rect 16 305 23 308
rect 25 318 33 327
rect 25 316 28 318
rect 30 316 33 318
rect 25 305 33 316
rect 35 325 43 327
rect 35 323 38 325
rect 40 323 43 325
rect 35 318 43 323
rect 35 316 38 318
rect 40 316 43 318
rect 35 311 43 316
rect 35 309 38 311
rect 40 309 43 311
rect 35 305 43 309
rect 45 325 57 327
rect 45 323 52 325
rect 54 323 57 325
rect 45 305 57 323
rect 59 317 64 327
rect 68 325 75 327
rect 68 323 70 325
rect 72 323 75 325
rect 68 321 75 323
rect 59 309 66 317
rect 70 314 75 321
rect 77 319 86 327
rect 107 320 112 327
rect 77 314 88 319
rect 79 309 88 314
rect 90 317 97 319
rect 90 315 93 317
rect 95 315 97 317
rect 90 313 97 315
rect 105 318 112 320
rect 105 316 107 318
rect 109 316 112 318
rect 105 314 112 316
rect 114 314 123 327
rect 90 309 95 313
rect 116 310 123 314
rect 59 307 62 309
rect 64 307 66 309
rect 59 305 66 307
rect 79 307 81 309
rect 83 307 86 309
rect 79 305 86 307
rect 116 308 118 310
rect 120 308 123 310
rect 116 305 123 308
rect 125 318 133 327
rect 125 316 128 318
rect 130 316 133 318
rect 125 305 133 316
rect 135 325 143 327
rect 135 323 138 325
rect 140 323 143 325
rect 135 318 143 323
rect 135 316 138 318
rect 140 316 143 318
rect 135 311 143 316
rect 135 309 138 311
rect 140 309 143 311
rect 135 305 143 309
rect 145 325 157 327
rect 145 323 152 325
rect 154 323 157 325
rect 145 305 157 323
rect 159 317 164 327
rect 168 325 175 327
rect 168 323 170 325
rect 172 323 175 325
rect 168 321 175 323
rect 159 309 166 317
rect 170 314 175 321
rect 177 319 186 327
rect 207 320 212 327
rect 177 314 188 319
rect 179 309 188 314
rect 190 317 197 319
rect 190 315 193 317
rect 195 315 197 317
rect 190 313 197 315
rect 205 318 212 320
rect 205 316 207 318
rect 209 316 212 318
rect 205 314 212 316
rect 214 314 223 327
rect 190 309 195 313
rect 216 310 223 314
rect 159 307 162 309
rect 164 307 166 309
rect 159 305 166 307
rect 179 307 181 309
rect 183 307 186 309
rect 179 305 186 307
rect 216 308 218 310
rect 220 308 223 310
rect 216 305 223 308
rect 225 318 233 327
rect 225 316 228 318
rect 230 316 233 318
rect 225 305 233 316
rect 235 325 243 327
rect 235 323 238 325
rect 240 323 243 325
rect 235 318 243 323
rect 235 316 238 318
rect 240 316 243 318
rect 235 311 243 316
rect 235 309 238 311
rect 240 309 243 311
rect 235 305 243 309
rect 245 325 257 327
rect 245 323 252 325
rect 254 323 257 325
rect 245 305 257 323
rect 259 317 264 327
rect 268 325 275 327
rect 268 323 270 325
rect 272 323 275 325
rect 268 321 275 323
rect 259 309 266 317
rect 270 314 275 321
rect 277 319 286 327
rect 307 320 312 327
rect 277 314 288 319
rect 279 309 288 314
rect 290 317 297 319
rect 290 315 293 317
rect 295 315 297 317
rect 290 313 297 315
rect 305 318 312 320
rect 305 316 307 318
rect 309 316 312 318
rect 305 314 312 316
rect 314 314 323 327
rect 290 309 295 313
rect 316 310 323 314
rect 259 307 262 309
rect 264 307 266 309
rect 259 305 266 307
rect 279 307 281 309
rect 283 307 286 309
rect 279 305 286 307
rect 316 308 318 310
rect 320 308 323 310
rect 316 305 323 308
rect 325 318 333 327
rect 325 316 328 318
rect 330 316 333 318
rect 325 305 333 316
rect 335 318 343 327
rect 335 316 338 318
rect 340 316 343 318
rect 335 311 343 316
rect 335 309 338 311
rect 340 309 343 311
rect 335 305 343 309
rect 345 325 357 327
rect 345 323 352 325
rect 354 323 357 325
rect 345 305 357 323
rect 359 317 364 327
rect 368 325 375 327
rect 368 323 370 325
rect 372 323 375 325
rect 368 321 375 323
rect 359 309 366 317
rect 370 314 375 321
rect 377 319 386 327
rect 407 320 412 327
rect 377 314 388 319
rect 379 309 388 314
rect 390 317 397 319
rect 390 315 393 317
rect 395 315 397 317
rect 390 313 397 315
rect 405 318 412 320
rect 405 316 407 318
rect 409 316 412 318
rect 405 314 412 316
rect 414 314 423 327
rect 390 309 395 313
rect 416 310 423 314
rect 359 307 362 309
rect 364 307 366 309
rect 359 305 366 307
rect 379 307 381 309
rect 383 307 386 309
rect 379 305 386 307
rect 416 308 418 310
rect 420 308 423 310
rect 416 305 423 308
rect 425 318 433 327
rect 425 316 428 318
rect 430 316 433 318
rect 425 305 433 316
rect 435 325 443 327
rect 435 323 438 325
rect 440 323 443 325
rect 435 318 443 323
rect 435 316 438 318
rect 440 316 443 318
rect 435 311 443 316
rect 435 309 438 311
rect 440 309 443 311
rect 435 305 443 309
rect 445 325 457 327
rect 445 323 452 325
rect 454 323 457 325
rect 445 305 457 323
rect 459 317 464 327
rect 468 325 475 327
rect 468 323 470 325
rect 472 323 475 325
rect 468 321 475 323
rect 459 309 466 317
rect 470 314 475 321
rect 477 319 486 327
rect 507 320 512 327
rect 477 314 488 319
rect 479 309 488 314
rect 490 317 497 319
rect 490 315 493 317
rect 495 315 497 317
rect 490 313 497 315
rect 505 318 512 320
rect 505 316 507 318
rect 509 316 512 318
rect 505 314 512 316
rect 514 314 523 327
rect 490 309 495 313
rect 516 310 523 314
rect 459 307 462 309
rect 464 307 466 309
rect 459 305 466 307
rect 479 307 481 309
rect 483 307 486 309
rect 479 305 486 307
rect 516 308 518 310
rect 520 308 523 310
rect 516 305 523 308
rect 525 318 533 327
rect 525 316 528 318
rect 530 316 533 318
rect 525 305 533 316
rect 535 325 543 327
rect 535 323 538 325
rect 540 323 543 325
rect 535 318 543 323
rect 535 316 538 318
rect 540 316 543 318
rect 535 311 543 316
rect 535 309 538 311
rect 540 309 543 311
rect 535 305 543 309
rect 545 325 557 327
rect 545 323 552 325
rect 554 323 557 325
rect 545 305 557 323
rect 559 317 564 327
rect 568 325 575 327
rect 568 323 570 325
rect 572 323 575 325
rect 568 321 575 323
rect 559 309 566 317
rect 570 314 575 321
rect 577 319 586 327
rect 607 320 612 327
rect 577 314 588 319
rect 579 309 588 314
rect 590 317 597 319
rect 590 315 593 317
rect 595 315 597 317
rect 590 313 597 315
rect 605 318 612 320
rect 605 316 607 318
rect 609 316 612 318
rect 605 314 612 316
rect 614 314 623 327
rect 590 309 595 313
rect 616 310 623 314
rect 559 307 562 309
rect 564 307 566 309
rect 559 305 566 307
rect 579 307 581 309
rect 583 307 586 309
rect 579 305 586 307
rect 616 308 618 310
rect 620 308 623 310
rect 616 305 623 308
rect 625 318 633 327
rect 625 316 628 318
rect 630 316 633 318
rect 625 305 633 316
rect 635 325 643 327
rect 635 323 638 325
rect 640 323 643 325
rect 635 318 643 323
rect 635 316 638 318
rect 640 316 643 318
rect 635 311 643 316
rect 635 309 638 311
rect 640 309 643 311
rect 635 305 643 309
rect 645 325 657 327
rect 645 323 652 325
rect 654 323 657 325
rect 645 305 657 323
rect 659 317 664 327
rect 668 325 675 327
rect 668 323 670 325
rect 672 323 675 325
rect 668 321 675 323
rect 659 309 666 317
rect 670 314 675 321
rect 677 319 686 327
rect 707 320 712 327
rect 677 314 688 319
rect 679 309 688 314
rect 690 317 697 319
rect 690 315 693 317
rect 695 315 697 317
rect 690 313 697 315
rect 705 318 712 320
rect 705 316 707 318
rect 709 316 712 318
rect 705 314 712 316
rect 714 314 723 327
rect 690 309 695 313
rect 716 310 723 314
rect 659 307 662 309
rect 664 307 666 309
rect 659 305 666 307
rect 679 307 681 309
rect 683 307 686 309
rect 679 305 686 307
rect 716 308 718 310
rect 720 308 723 310
rect 716 305 723 308
rect 725 318 733 327
rect 725 316 728 318
rect 730 316 733 318
rect 725 305 733 316
rect 735 325 743 327
rect 735 323 738 325
rect 740 323 743 325
rect 735 318 743 323
rect 735 316 738 318
rect 740 316 743 318
rect 735 311 743 316
rect 735 309 738 311
rect 740 309 743 311
rect 735 305 743 309
rect 745 325 757 327
rect 745 323 752 325
rect 754 323 757 325
rect 745 305 757 323
rect 759 317 764 327
rect 768 325 775 327
rect 768 323 770 325
rect 772 323 775 325
rect 768 321 775 323
rect 759 309 766 317
rect 770 314 775 321
rect 777 319 786 327
rect 777 314 788 319
rect 779 309 788 314
rect 790 317 797 319
rect 790 315 793 317
rect 795 315 797 317
rect 790 313 797 315
rect 790 309 795 313
rect 759 307 762 309
rect 764 307 766 309
rect 759 305 766 307
rect 779 307 781 309
rect 783 307 786 309
rect 779 305 786 307
rect 16 279 23 281
rect 16 277 19 279
rect 21 277 23 279
rect 36 279 43 281
rect 36 277 38 279
rect 40 277 43 279
rect 7 273 12 277
rect 5 271 12 273
rect 5 269 7 271
rect 9 269 12 271
rect 5 267 12 269
rect 14 272 23 277
rect 14 267 25 272
rect 16 259 25 267
rect 27 265 32 272
rect 36 269 43 277
rect 27 263 34 265
rect 27 261 30 263
rect 32 261 34 263
rect 27 259 34 261
rect 38 259 43 269
rect 45 263 57 281
rect 45 261 48 263
rect 50 261 57 263
rect 45 259 57 261
rect 59 277 67 281
rect 59 275 62 277
rect 64 275 67 277
rect 59 270 67 275
rect 59 268 62 270
rect 64 268 67 270
rect 59 263 67 268
rect 59 261 62 263
rect 64 261 67 263
rect 59 259 67 261
rect 69 270 77 281
rect 69 268 72 270
rect 74 268 77 270
rect 69 259 77 268
rect 79 278 86 281
rect 79 276 82 278
rect 84 276 86 278
rect 116 279 123 281
rect 116 277 119 279
rect 121 277 123 279
rect 136 279 143 281
rect 136 277 138 279
rect 140 277 143 279
rect 79 272 86 276
rect 107 273 112 277
rect 79 259 88 272
rect 90 270 97 272
rect 90 268 93 270
rect 95 268 97 270
rect 90 266 97 268
rect 105 271 112 273
rect 105 269 107 271
rect 109 269 112 271
rect 105 267 112 269
rect 114 272 123 277
rect 114 267 125 272
rect 90 259 95 266
rect 116 259 125 267
rect 127 265 132 272
rect 136 269 143 277
rect 127 263 134 265
rect 127 261 130 263
rect 132 261 134 263
rect 127 259 134 261
rect 138 259 143 269
rect 145 263 157 281
rect 145 261 148 263
rect 150 261 157 263
rect 145 259 157 261
rect 159 277 167 281
rect 159 275 162 277
rect 164 275 167 277
rect 159 270 167 275
rect 159 268 162 270
rect 164 268 167 270
rect 159 263 167 268
rect 159 261 162 263
rect 164 261 167 263
rect 159 259 167 261
rect 169 270 177 281
rect 169 268 172 270
rect 174 268 177 270
rect 169 259 177 268
rect 179 278 186 281
rect 179 276 182 278
rect 184 276 186 278
rect 216 279 223 281
rect 216 277 219 279
rect 221 277 223 279
rect 236 279 243 281
rect 236 277 238 279
rect 240 277 243 279
rect 179 272 186 276
rect 207 273 212 277
rect 179 259 188 272
rect 190 270 197 272
rect 190 268 193 270
rect 195 268 197 270
rect 190 266 197 268
rect 205 271 212 273
rect 205 269 207 271
rect 209 269 212 271
rect 205 267 212 269
rect 214 272 223 277
rect 214 267 225 272
rect 190 259 195 266
rect 216 259 225 267
rect 227 265 232 272
rect 236 269 243 277
rect 227 263 234 265
rect 227 261 230 263
rect 232 261 234 263
rect 227 259 234 261
rect 238 259 243 269
rect 245 263 257 281
rect 245 261 248 263
rect 250 261 257 263
rect 245 259 257 261
rect 259 277 267 281
rect 259 275 262 277
rect 264 275 267 277
rect 259 270 267 275
rect 259 268 262 270
rect 264 268 267 270
rect 259 263 267 268
rect 259 261 262 263
rect 264 261 267 263
rect 259 259 267 261
rect 269 270 277 281
rect 269 268 272 270
rect 274 268 277 270
rect 269 259 277 268
rect 279 278 286 281
rect 279 276 282 278
rect 284 276 286 278
rect 316 279 323 281
rect 316 277 319 279
rect 321 277 323 279
rect 336 279 343 281
rect 336 277 338 279
rect 340 277 343 279
rect 279 273 286 276
rect 307 273 312 277
rect 279 259 288 273
rect 290 271 297 273
rect 290 269 293 271
rect 295 269 297 271
rect 290 266 297 269
rect 305 271 312 273
rect 305 269 307 271
rect 309 269 312 271
rect 305 267 312 269
rect 314 272 323 277
rect 314 267 325 272
rect 290 259 295 266
rect 316 259 325 267
rect 327 265 332 272
rect 336 269 343 277
rect 327 263 334 265
rect 327 261 330 263
rect 332 261 334 263
rect 327 259 334 261
rect 338 259 343 269
rect 345 263 357 281
rect 345 261 348 263
rect 350 261 357 263
rect 345 259 357 261
rect 359 277 367 281
rect 359 275 362 277
rect 364 275 367 277
rect 359 270 367 275
rect 359 268 362 270
rect 364 268 367 270
rect 359 263 367 268
rect 359 261 362 263
rect 364 261 367 263
rect 359 259 367 261
rect 369 270 377 281
rect 369 268 372 270
rect 374 268 377 270
rect 369 259 377 268
rect 379 278 386 281
rect 379 276 382 278
rect 384 276 386 278
rect 418 279 425 281
rect 418 277 421 279
rect 423 277 425 279
rect 438 279 445 281
rect 438 277 440 279
rect 442 277 445 279
rect 379 272 386 276
rect 409 273 414 277
rect 379 259 388 272
rect 390 270 397 272
rect 390 268 393 270
rect 395 268 397 270
rect 390 266 397 268
rect 407 271 414 273
rect 407 269 409 271
rect 411 269 414 271
rect 407 267 414 269
rect 416 272 425 277
rect 416 267 427 272
rect 390 259 395 266
rect 418 259 427 267
rect 429 265 434 272
rect 438 269 445 277
rect 429 263 436 265
rect 429 261 432 263
rect 434 261 436 263
rect 429 259 436 261
rect 440 259 445 269
rect 447 263 459 281
rect 447 261 450 263
rect 452 261 459 263
rect 447 259 459 261
rect 461 277 469 281
rect 461 275 464 277
rect 466 275 469 277
rect 461 270 469 275
rect 461 268 464 270
rect 466 268 469 270
rect 461 263 469 268
rect 461 261 464 263
rect 466 261 469 263
rect 461 259 469 261
rect 471 270 479 281
rect 471 268 474 270
rect 476 268 479 270
rect 471 259 479 268
rect 481 278 488 281
rect 481 276 484 278
rect 486 276 488 278
rect 518 279 525 281
rect 518 277 521 279
rect 523 277 525 279
rect 538 279 545 281
rect 538 277 540 279
rect 542 277 545 279
rect 481 273 488 276
rect 509 273 514 277
rect 481 260 490 273
rect 492 271 499 273
rect 492 269 495 271
rect 497 269 499 271
rect 492 266 499 269
rect 507 271 514 273
rect 507 269 509 271
rect 511 269 514 271
rect 507 267 514 269
rect 516 272 525 277
rect 516 267 527 272
rect 492 260 497 266
rect 481 259 488 260
rect 518 259 527 267
rect 529 265 534 272
rect 538 269 545 277
rect 529 263 536 265
rect 529 261 532 263
rect 534 261 536 263
rect 529 259 536 261
rect 540 259 545 269
rect 547 263 559 281
rect 547 261 550 263
rect 552 261 559 263
rect 547 259 559 261
rect 561 277 569 281
rect 561 275 564 277
rect 566 275 569 277
rect 561 270 569 275
rect 561 268 564 270
rect 566 268 569 270
rect 561 263 569 268
rect 561 261 564 263
rect 566 261 569 263
rect 561 259 569 261
rect 571 270 579 281
rect 571 268 574 270
rect 576 268 579 270
rect 571 259 579 268
rect 581 278 588 281
rect 581 276 584 278
rect 586 276 588 278
rect 618 279 625 281
rect 618 277 621 279
rect 623 277 625 279
rect 638 279 645 281
rect 638 277 640 279
rect 642 277 645 279
rect 581 272 588 276
rect 609 273 614 277
rect 581 259 590 272
rect 592 270 599 272
rect 592 268 595 270
rect 597 268 599 270
rect 592 266 599 268
rect 607 271 614 273
rect 607 269 609 271
rect 611 269 614 271
rect 607 267 614 269
rect 616 272 625 277
rect 616 267 627 272
rect 592 259 597 266
rect 618 259 627 267
rect 629 265 634 272
rect 638 269 645 277
rect 629 263 636 265
rect 629 261 632 263
rect 634 261 636 263
rect 629 259 636 261
rect 640 259 645 269
rect 647 263 659 281
rect 647 261 650 263
rect 652 261 659 263
rect 647 259 659 261
rect 661 277 669 281
rect 661 275 664 277
rect 666 275 669 277
rect 661 270 669 275
rect 661 268 664 270
rect 666 268 669 270
rect 661 263 669 268
rect 661 261 664 263
rect 666 261 669 263
rect 661 259 669 261
rect 671 270 679 281
rect 671 268 674 270
rect 676 268 679 270
rect 671 259 679 268
rect 681 278 688 281
rect 681 276 684 278
rect 686 276 688 278
rect 718 279 725 281
rect 718 277 721 279
rect 723 277 725 279
rect 738 279 745 281
rect 738 277 740 279
rect 742 277 745 279
rect 681 273 688 276
rect 709 273 714 277
rect 681 260 690 273
rect 692 271 699 273
rect 692 269 695 271
rect 697 269 699 271
rect 692 266 699 269
rect 707 271 714 273
rect 707 269 709 271
rect 711 269 714 271
rect 707 267 714 269
rect 716 272 725 277
rect 716 267 727 272
rect 692 260 697 266
rect 681 259 688 260
rect 718 259 727 267
rect 729 265 734 272
rect 738 269 745 277
rect 729 263 736 265
rect 729 261 732 263
rect 734 261 736 263
rect 729 259 736 261
rect 740 259 745 269
rect 747 263 759 281
rect 747 261 750 263
rect 752 261 759 263
rect 747 259 759 261
rect 761 277 769 281
rect 761 275 764 277
rect 766 275 769 277
rect 761 270 769 275
rect 761 268 764 270
rect 766 268 769 270
rect 761 263 769 268
rect 761 261 764 263
rect 766 261 769 263
rect 761 259 769 261
rect 771 270 779 281
rect 771 268 774 270
rect 776 268 779 270
rect 771 259 779 268
rect 781 278 788 281
rect 781 276 784 278
rect 786 276 788 278
rect 781 272 788 276
rect 781 259 790 272
rect 792 270 799 272
rect 792 268 795 270
rect 797 268 799 270
rect 792 266 799 268
rect 792 259 797 266
rect 16 175 25 183
rect 5 173 12 175
rect 5 171 7 173
rect 9 171 12 173
rect 5 169 12 171
rect 7 165 12 169
rect 14 170 25 175
rect 27 181 34 183
rect 27 179 30 181
rect 32 179 34 181
rect 27 177 34 179
rect 27 170 32 177
rect 38 173 43 183
rect 14 165 23 170
rect 36 165 43 173
rect 16 163 19 165
rect 21 163 23 165
rect 16 161 23 163
rect 36 163 38 165
rect 40 163 43 165
rect 36 161 43 163
rect 45 181 57 183
rect 45 179 48 181
rect 50 179 57 181
rect 45 161 57 179
rect 59 181 67 183
rect 59 179 62 181
rect 64 179 67 181
rect 59 174 67 179
rect 59 172 62 174
rect 64 172 67 174
rect 59 167 67 172
rect 59 165 62 167
rect 64 165 67 167
rect 59 161 67 165
rect 69 174 77 183
rect 69 172 72 174
rect 74 172 77 174
rect 69 161 77 172
rect 79 170 88 183
rect 90 176 95 183
rect 90 174 97 176
rect 116 175 125 183
rect 90 172 93 174
rect 95 172 97 174
rect 90 170 97 172
rect 105 173 112 175
rect 105 171 107 173
rect 109 171 112 173
rect 79 166 86 170
rect 79 164 82 166
rect 84 164 86 166
rect 105 169 112 171
rect 107 165 112 169
rect 114 170 125 175
rect 127 181 134 183
rect 127 179 130 181
rect 132 179 134 181
rect 127 177 134 179
rect 127 170 132 177
rect 138 173 143 183
rect 114 165 123 170
rect 136 165 143 173
rect 79 161 86 164
rect 116 163 119 165
rect 121 163 123 165
rect 116 161 123 163
rect 136 163 138 165
rect 140 163 143 165
rect 136 161 143 163
rect 145 181 157 183
rect 145 179 148 181
rect 150 179 157 181
rect 145 161 157 179
rect 159 181 167 183
rect 159 179 162 181
rect 164 179 167 181
rect 159 174 167 179
rect 159 172 162 174
rect 164 172 167 174
rect 159 167 167 172
rect 159 165 162 167
rect 164 165 167 167
rect 159 161 167 165
rect 169 174 177 183
rect 169 172 172 174
rect 174 172 177 174
rect 169 161 177 172
rect 179 170 188 183
rect 190 176 195 183
rect 190 174 197 176
rect 216 175 225 183
rect 190 172 193 174
rect 195 172 197 174
rect 190 170 197 172
rect 205 173 212 175
rect 205 171 207 173
rect 209 171 212 173
rect 179 166 186 170
rect 179 164 182 166
rect 184 164 186 166
rect 205 169 212 171
rect 207 165 212 169
rect 214 170 225 175
rect 227 181 234 183
rect 227 179 230 181
rect 232 179 234 181
rect 227 177 234 179
rect 227 170 232 177
rect 238 173 243 183
rect 214 165 223 170
rect 236 165 243 173
rect 179 161 186 164
rect 216 163 219 165
rect 221 163 223 165
rect 216 161 223 163
rect 236 163 238 165
rect 240 163 243 165
rect 236 161 243 163
rect 245 181 257 183
rect 245 179 248 181
rect 250 179 257 181
rect 245 161 257 179
rect 259 181 267 183
rect 259 179 262 181
rect 264 179 267 181
rect 259 174 267 179
rect 259 172 262 174
rect 264 172 267 174
rect 259 167 267 172
rect 259 165 262 167
rect 264 165 267 167
rect 259 161 267 165
rect 269 174 277 183
rect 269 172 272 174
rect 274 172 277 174
rect 269 161 277 172
rect 279 170 288 183
rect 290 176 295 183
rect 290 174 297 176
rect 316 175 325 183
rect 290 172 293 174
rect 295 172 297 174
rect 290 170 297 172
rect 305 173 312 175
rect 305 171 307 173
rect 309 171 312 173
rect 279 166 286 170
rect 279 164 282 166
rect 284 164 286 166
rect 305 169 312 171
rect 307 165 312 169
rect 314 170 325 175
rect 327 181 334 183
rect 327 179 330 181
rect 332 179 334 181
rect 327 177 334 179
rect 327 170 332 177
rect 338 173 343 183
rect 314 165 323 170
rect 336 165 343 173
rect 279 161 286 164
rect 316 163 319 165
rect 321 163 323 165
rect 316 161 323 163
rect 336 163 338 165
rect 340 163 343 165
rect 336 161 343 163
rect 345 181 357 183
rect 345 179 348 181
rect 350 179 357 181
rect 345 161 357 179
rect 359 181 367 183
rect 359 179 362 181
rect 364 179 367 181
rect 359 174 367 179
rect 359 172 362 174
rect 364 172 367 174
rect 359 167 367 172
rect 359 165 362 167
rect 364 165 367 167
rect 359 161 367 165
rect 369 174 377 183
rect 369 172 372 174
rect 374 172 377 174
rect 369 161 377 172
rect 379 170 388 183
rect 390 176 395 183
rect 390 174 397 176
rect 418 175 427 183
rect 390 172 393 174
rect 395 172 397 174
rect 390 170 397 172
rect 407 173 414 175
rect 407 171 409 173
rect 411 171 414 173
rect 379 166 386 170
rect 379 164 382 166
rect 384 164 386 166
rect 407 169 414 171
rect 409 165 414 169
rect 416 170 427 175
rect 429 181 436 183
rect 429 179 432 181
rect 434 179 436 181
rect 429 177 436 179
rect 429 170 434 177
rect 440 173 445 183
rect 416 165 425 170
rect 438 165 445 173
rect 379 161 386 164
rect 418 163 421 165
rect 423 163 425 165
rect 418 161 425 163
rect 438 163 440 165
rect 442 163 445 165
rect 438 161 445 163
rect 447 181 459 183
rect 447 179 450 181
rect 452 179 459 181
rect 447 161 459 179
rect 461 181 469 183
rect 461 179 464 181
rect 466 179 469 181
rect 461 174 469 179
rect 461 172 464 174
rect 466 172 469 174
rect 461 167 469 172
rect 461 165 464 167
rect 466 165 469 167
rect 461 161 469 165
rect 471 174 479 183
rect 471 172 474 174
rect 476 172 479 174
rect 471 161 479 172
rect 481 170 490 183
rect 492 176 497 183
rect 492 174 499 176
rect 518 175 527 183
rect 492 172 495 174
rect 497 172 499 174
rect 492 170 499 172
rect 507 173 514 175
rect 507 171 509 173
rect 511 171 514 173
rect 481 166 488 170
rect 481 164 484 166
rect 486 164 488 166
rect 507 169 514 171
rect 509 165 514 169
rect 516 170 527 175
rect 529 181 536 183
rect 529 179 532 181
rect 534 179 536 181
rect 529 177 536 179
rect 529 170 534 177
rect 540 173 545 183
rect 516 165 525 170
rect 538 165 545 173
rect 481 161 488 164
rect 518 163 521 165
rect 523 163 525 165
rect 518 161 525 163
rect 538 163 540 165
rect 542 163 545 165
rect 538 161 545 163
rect 547 181 559 183
rect 547 179 550 181
rect 552 179 559 181
rect 547 161 559 179
rect 561 181 569 183
rect 561 179 564 181
rect 566 179 569 181
rect 561 174 569 179
rect 561 172 564 174
rect 566 172 569 174
rect 561 167 569 172
rect 561 165 564 167
rect 566 165 569 167
rect 561 161 569 165
rect 571 174 579 183
rect 571 172 574 174
rect 576 172 579 174
rect 571 161 579 172
rect 581 170 590 183
rect 592 176 597 183
rect 592 174 599 176
rect 618 175 627 183
rect 592 172 595 174
rect 597 172 599 174
rect 592 170 599 172
rect 607 173 614 175
rect 607 171 609 173
rect 611 171 614 173
rect 581 166 588 170
rect 581 164 584 166
rect 586 164 588 166
rect 607 169 614 171
rect 609 165 614 169
rect 616 170 627 175
rect 629 181 636 183
rect 629 179 632 181
rect 634 179 636 181
rect 629 177 636 179
rect 629 170 634 177
rect 640 173 645 183
rect 616 165 625 170
rect 638 165 645 173
rect 581 161 588 164
rect 618 163 621 165
rect 623 163 625 165
rect 618 161 625 163
rect 638 163 640 165
rect 642 163 645 165
rect 638 161 645 163
rect 647 181 659 183
rect 647 179 650 181
rect 652 179 659 181
rect 647 161 659 179
rect 661 181 669 183
rect 661 179 664 181
rect 666 179 669 181
rect 661 174 669 179
rect 661 172 664 174
rect 666 172 669 174
rect 661 167 669 172
rect 661 165 664 167
rect 666 165 669 167
rect 661 161 669 165
rect 671 174 679 183
rect 671 172 674 174
rect 676 172 679 174
rect 671 161 679 172
rect 681 170 690 183
rect 692 176 697 183
rect 692 174 699 176
rect 718 175 727 183
rect 692 172 695 174
rect 697 172 699 174
rect 692 170 699 172
rect 707 173 714 175
rect 707 171 709 173
rect 711 171 714 173
rect 681 166 688 170
rect 681 164 684 166
rect 686 164 688 166
rect 707 169 714 171
rect 709 165 714 169
rect 716 170 727 175
rect 729 181 736 183
rect 729 179 732 181
rect 734 179 736 181
rect 729 177 736 179
rect 729 170 734 177
rect 740 173 745 183
rect 716 165 725 170
rect 738 165 745 173
rect 681 161 688 164
rect 718 163 721 165
rect 723 163 725 165
rect 718 161 725 163
rect 738 163 740 165
rect 742 163 745 165
rect 738 161 745 163
rect 747 181 759 183
rect 747 179 750 181
rect 752 179 759 181
rect 747 161 759 179
rect 761 181 769 183
rect 761 179 764 181
rect 766 179 769 181
rect 761 174 769 179
rect 761 172 764 174
rect 766 172 769 174
rect 761 167 769 172
rect 761 165 764 167
rect 766 165 769 167
rect 761 161 769 165
rect 771 174 779 183
rect 771 172 774 174
rect 776 172 779 174
rect 771 161 779 172
rect 781 170 790 183
rect 792 176 797 183
rect 792 174 799 176
rect 792 172 795 174
rect 797 172 799 174
rect 792 170 799 172
rect 781 166 788 170
rect 781 164 784 166
rect 786 164 788 166
rect 781 161 788 164
rect 16 135 23 137
rect 16 133 19 135
rect 21 133 23 135
rect 36 135 43 137
rect 36 133 38 135
rect 40 133 43 135
rect 7 129 12 133
rect 5 127 12 129
rect 5 125 7 127
rect 9 125 12 127
rect 5 123 12 125
rect 14 128 23 133
rect 14 123 25 128
rect 16 115 25 123
rect 27 121 32 128
rect 36 125 43 133
rect 27 119 34 121
rect 27 117 30 119
rect 32 117 34 119
rect 27 115 34 117
rect 38 115 43 125
rect 45 119 57 137
rect 45 117 48 119
rect 50 117 57 119
rect 45 115 57 117
rect 59 133 67 137
rect 59 131 62 133
rect 64 131 67 133
rect 59 126 67 131
rect 59 124 62 126
rect 64 124 67 126
rect 59 119 67 124
rect 59 117 62 119
rect 64 117 67 119
rect 59 115 67 117
rect 69 126 77 137
rect 69 124 72 126
rect 74 124 77 126
rect 69 115 77 124
rect 79 134 86 137
rect 79 132 82 134
rect 84 132 86 134
rect 116 135 123 137
rect 116 133 119 135
rect 121 133 123 135
rect 136 135 143 137
rect 136 133 138 135
rect 140 133 143 135
rect 79 128 86 132
rect 107 129 112 133
rect 79 115 88 128
rect 90 126 97 128
rect 90 124 93 126
rect 95 124 97 126
rect 90 122 97 124
rect 105 127 112 129
rect 105 125 107 127
rect 109 125 112 127
rect 105 123 112 125
rect 114 128 123 133
rect 114 123 125 128
rect 90 115 95 122
rect 116 115 125 123
rect 127 121 132 128
rect 136 125 143 133
rect 127 119 134 121
rect 127 117 130 119
rect 132 117 134 119
rect 127 115 134 117
rect 138 115 143 125
rect 145 119 157 137
rect 145 117 148 119
rect 150 117 157 119
rect 145 115 157 117
rect 159 133 167 137
rect 159 131 162 133
rect 164 131 167 133
rect 159 126 167 131
rect 159 124 162 126
rect 164 124 167 126
rect 159 119 167 124
rect 159 117 162 119
rect 164 117 167 119
rect 159 115 167 117
rect 169 126 177 137
rect 169 124 172 126
rect 174 124 177 126
rect 169 115 177 124
rect 179 134 186 137
rect 179 132 182 134
rect 184 132 186 134
rect 216 135 223 137
rect 216 133 219 135
rect 221 133 223 135
rect 236 135 243 137
rect 236 133 238 135
rect 240 133 243 135
rect 179 128 186 132
rect 207 129 212 133
rect 179 115 188 128
rect 190 126 197 128
rect 190 124 193 126
rect 195 124 197 126
rect 190 122 197 124
rect 205 127 212 129
rect 205 125 207 127
rect 209 125 212 127
rect 205 123 212 125
rect 214 128 223 133
rect 214 123 225 128
rect 190 115 195 122
rect 216 115 225 123
rect 227 121 232 128
rect 236 125 243 133
rect 227 119 234 121
rect 227 117 230 119
rect 232 117 234 119
rect 227 115 234 117
rect 238 115 243 125
rect 245 119 257 137
rect 245 117 248 119
rect 250 117 257 119
rect 245 115 257 117
rect 259 133 267 137
rect 259 131 262 133
rect 264 131 267 133
rect 259 126 267 131
rect 259 124 262 126
rect 264 124 267 126
rect 259 119 267 124
rect 259 117 262 119
rect 264 117 267 119
rect 259 115 267 117
rect 269 126 277 137
rect 269 124 272 126
rect 274 124 277 126
rect 269 115 277 124
rect 279 134 286 137
rect 279 132 282 134
rect 284 132 286 134
rect 316 135 323 137
rect 316 133 319 135
rect 321 133 323 135
rect 336 135 343 137
rect 336 133 338 135
rect 340 133 343 135
rect 279 128 286 132
rect 307 129 312 133
rect 279 115 288 128
rect 290 126 297 128
rect 290 124 293 126
rect 295 124 297 126
rect 290 122 297 124
rect 305 127 312 129
rect 305 125 307 127
rect 309 125 312 127
rect 305 123 312 125
rect 314 128 323 133
rect 314 123 325 128
rect 290 115 295 122
rect 316 115 325 123
rect 327 121 332 128
rect 336 125 343 133
rect 327 119 334 121
rect 327 117 330 119
rect 332 117 334 119
rect 327 115 334 117
rect 338 115 343 125
rect 345 119 357 137
rect 345 117 348 119
rect 350 117 357 119
rect 345 115 357 117
rect 359 133 367 137
rect 359 131 362 133
rect 364 131 367 133
rect 359 126 367 131
rect 359 124 362 126
rect 364 124 367 126
rect 359 119 367 124
rect 359 117 362 119
rect 364 117 367 119
rect 359 115 367 117
rect 369 126 377 137
rect 369 124 372 126
rect 374 124 377 126
rect 369 115 377 124
rect 379 134 386 137
rect 379 132 382 134
rect 384 132 386 134
rect 418 135 425 137
rect 418 133 421 135
rect 423 133 425 135
rect 438 135 445 137
rect 438 133 440 135
rect 442 133 445 135
rect 379 128 386 132
rect 409 129 414 133
rect 379 115 388 128
rect 390 126 397 128
rect 390 124 393 126
rect 395 124 397 126
rect 390 122 397 124
rect 407 127 414 129
rect 407 125 409 127
rect 411 125 414 127
rect 407 123 414 125
rect 416 128 425 133
rect 416 123 427 128
rect 390 115 395 122
rect 418 115 427 123
rect 429 121 434 128
rect 438 125 445 133
rect 429 119 436 121
rect 429 117 432 119
rect 434 117 436 119
rect 429 115 436 117
rect 440 115 445 125
rect 447 119 459 137
rect 447 117 450 119
rect 452 117 459 119
rect 447 115 459 117
rect 461 133 469 137
rect 461 131 464 133
rect 466 131 469 133
rect 461 126 469 131
rect 461 124 464 126
rect 466 124 469 126
rect 461 119 469 124
rect 461 117 464 119
rect 466 117 469 119
rect 461 115 469 117
rect 471 126 479 137
rect 471 124 474 126
rect 476 124 479 126
rect 471 115 479 124
rect 481 134 488 137
rect 481 132 484 134
rect 486 132 488 134
rect 518 135 525 137
rect 518 133 521 135
rect 523 133 525 135
rect 538 135 545 137
rect 538 133 540 135
rect 542 133 545 135
rect 481 128 488 132
rect 509 129 514 133
rect 481 115 490 128
rect 492 126 499 128
rect 492 124 495 126
rect 497 124 499 126
rect 492 122 499 124
rect 507 127 514 129
rect 507 125 509 127
rect 511 125 514 127
rect 507 123 514 125
rect 516 128 525 133
rect 516 123 527 128
rect 492 115 497 122
rect 518 115 527 123
rect 529 121 534 128
rect 538 125 545 133
rect 529 119 536 121
rect 529 117 532 119
rect 534 117 536 119
rect 529 115 536 117
rect 540 115 545 125
rect 547 119 559 137
rect 547 117 550 119
rect 552 117 559 119
rect 547 115 559 117
rect 561 133 569 137
rect 561 131 564 133
rect 566 131 569 133
rect 561 126 569 131
rect 561 124 564 126
rect 566 124 569 126
rect 561 119 569 124
rect 561 117 564 119
rect 566 117 569 119
rect 561 115 569 117
rect 571 126 579 137
rect 571 124 574 126
rect 576 124 579 126
rect 571 115 579 124
rect 581 134 588 137
rect 581 132 584 134
rect 586 132 588 134
rect 618 135 625 137
rect 618 133 621 135
rect 623 133 625 135
rect 638 135 645 137
rect 638 133 640 135
rect 642 133 645 135
rect 581 128 588 132
rect 609 129 614 133
rect 581 115 590 128
rect 592 126 599 128
rect 592 124 595 126
rect 597 124 599 126
rect 592 122 599 124
rect 607 127 614 129
rect 607 125 609 127
rect 611 125 614 127
rect 607 123 614 125
rect 616 128 625 133
rect 616 123 627 128
rect 592 115 597 122
rect 618 115 627 123
rect 629 121 634 128
rect 638 125 645 133
rect 629 119 636 121
rect 629 117 632 119
rect 634 117 636 119
rect 629 115 636 117
rect 640 115 645 125
rect 647 119 659 137
rect 647 117 650 119
rect 652 117 659 119
rect 647 115 659 117
rect 661 133 669 137
rect 661 131 664 133
rect 666 131 669 133
rect 661 126 669 131
rect 661 124 664 126
rect 666 124 669 126
rect 661 119 669 124
rect 661 117 664 119
rect 666 117 669 119
rect 661 115 669 117
rect 671 126 679 137
rect 671 124 674 126
rect 676 124 679 126
rect 671 115 679 124
rect 681 134 688 137
rect 681 132 684 134
rect 686 132 688 134
rect 718 135 725 137
rect 718 133 721 135
rect 723 133 725 135
rect 738 135 745 137
rect 738 133 740 135
rect 742 133 745 135
rect 681 128 688 132
rect 709 129 714 133
rect 681 115 690 128
rect 692 126 699 128
rect 692 124 695 126
rect 697 124 699 126
rect 692 122 699 124
rect 707 127 714 129
rect 707 125 709 127
rect 711 125 714 127
rect 707 123 714 125
rect 716 128 725 133
rect 716 123 727 128
rect 692 115 697 122
rect 718 115 727 123
rect 729 121 734 128
rect 738 125 745 133
rect 729 119 736 121
rect 729 117 732 119
rect 734 117 736 119
rect 729 115 736 117
rect 740 115 745 125
rect 747 119 759 137
rect 747 117 750 119
rect 752 117 759 119
rect 747 115 759 117
rect 761 133 769 137
rect 761 131 764 133
rect 766 131 769 133
rect 761 126 769 131
rect 761 124 764 126
rect 766 124 769 126
rect 761 119 769 124
rect 761 117 764 119
rect 766 117 769 119
rect 761 115 769 117
rect 771 126 779 137
rect 771 124 774 126
rect 776 124 779 126
rect 771 115 779 124
rect 781 134 788 137
rect 781 132 784 134
rect 786 132 788 134
rect 781 128 788 132
rect 781 115 790 128
rect 792 126 799 128
rect 792 124 795 126
rect 797 124 799 126
rect 792 122 799 124
rect 792 115 797 122
rect 7 32 12 39
rect 5 30 12 32
rect 5 28 7 30
rect 9 28 12 30
rect 5 26 12 28
rect 14 26 23 39
rect 16 22 23 26
rect 16 20 18 22
rect 20 20 23 22
rect 16 17 23 20
rect 25 30 33 39
rect 25 28 28 30
rect 30 28 33 30
rect 25 17 33 28
rect 35 37 43 39
rect 35 35 38 37
rect 40 35 43 37
rect 35 30 43 35
rect 35 28 38 30
rect 40 28 43 30
rect 35 23 43 28
rect 35 21 38 23
rect 40 21 43 23
rect 35 17 43 21
rect 45 37 57 39
rect 45 35 52 37
rect 54 35 57 37
rect 45 17 57 35
rect 59 29 64 39
rect 68 37 75 39
rect 68 35 70 37
rect 72 35 75 37
rect 68 33 75 35
rect 59 21 66 29
rect 70 26 75 33
rect 77 31 86 39
rect 107 32 112 39
rect 77 26 88 31
rect 79 21 88 26
rect 90 29 97 31
rect 90 27 93 29
rect 95 27 97 29
rect 90 25 97 27
rect 105 30 112 32
rect 105 28 107 30
rect 109 28 112 30
rect 105 26 112 28
rect 114 26 123 39
rect 90 21 95 25
rect 116 22 123 26
rect 59 19 62 21
rect 64 19 66 21
rect 59 17 66 19
rect 79 19 81 21
rect 83 19 86 21
rect 79 17 86 19
rect 116 20 118 22
rect 120 20 123 22
rect 116 17 123 20
rect 125 30 133 39
rect 125 28 128 30
rect 130 28 133 30
rect 125 17 133 28
rect 135 37 143 39
rect 135 35 138 37
rect 140 35 143 37
rect 135 30 143 35
rect 135 28 138 30
rect 140 28 143 30
rect 135 23 143 28
rect 135 21 138 23
rect 140 21 143 23
rect 135 17 143 21
rect 145 37 157 39
rect 145 35 152 37
rect 154 35 157 37
rect 145 17 157 35
rect 159 29 164 39
rect 168 37 175 39
rect 168 35 170 37
rect 172 35 175 37
rect 168 33 175 35
rect 159 21 166 29
rect 170 26 175 33
rect 177 31 186 39
rect 207 32 212 39
rect 177 26 188 31
rect 179 21 188 26
rect 190 29 197 31
rect 190 27 193 29
rect 195 27 197 29
rect 190 25 197 27
rect 205 30 212 32
rect 205 28 207 30
rect 209 28 212 30
rect 205 26 212 28
rect 214 26 223 39
rect 190 21 195 25
rect 216 22 223 26
rect 159 19 162 21
rect 164 19 166 21
rect 159 17 166 19
rect 179 19 181 21
rect 183 19 186 21
rect 179 17 186 19
rect 216 20 218 22
rect 220 20 223 22
rect 216 17 223 20
rect 225 30 233 39
rect 225 28 228 30
rect 230 28 233 30
rect 225 17 233 28
rect 235 37 243 39
rect 235 35 238 37
rect 240 35 243 37
rect 235 30 243 35
rect 235 28 238 30
rect 240 28 243 30
rect 235 23 243 28
rect 235 21 238 23
rect 240 21 243 23
rect 235 17 243 21
rect 245 37 257 39
rect 245 35 252 37
rect 254 35 257 37
rect 245 17 257 35
rect 259 29 264 39
rect 268 37 275 39
rect 268 35 270 37
rect 272 35 275 37
rect 268 33 275 35
rect 259 21 266 29
rect 270 26 275 33
rect 277 31 286 39
rect 307 32 312 39
rect 277 26 288 31
rect 279 21 288 26
rect 290 29 297 31
rect 290 27 293 29
rect 295 27 297 29
rect 290 25 297 27
rect 305 30 312 32
rect 305 28 307 30
rect 309 28 312 30
rect 305 26 312 28
rect 314 26 323 39
rect 290 21 295 25
rect 316 22 323 26
rect 259 19 262 21
rect 264 19 266 21
rect 259 17 266 19
rect 279 19 281 21
rect 283 19 286 21
rect 279 17 286 19
rect 316 20 318 22
rect 320 20 323 22
rect 316 17 323 20
rect 325 30 333 39
rect 325 28 328 30
rect 330 28 333 30
rect 325 17 333 28
rect 335 37 343 39
rect 335 35 338 37
rect 340 35 343 37
rect 335 30 343 35
rect 335 28 338 30
rect 340 28 343 30
rect 335 23 343 28
rect 335 21 338 23
rect 340 21 343 23
rect 335 17 343 21
rect 345 37 357 39
rect 345 35 352 37
rect 354 35 357 37
rect 345 17 357 35
rect 359 29 364 39
rect 368 37 375 39
rect 368 35 370 37
rect 372 35 375 37
rect 368 33 375 35
rect 359 21 366 29
rect 370 26 375 33
rect 377 31 386 39
rect 407 32 412 39
rect 377 26 388 31
rect 379 21 388 26
rect 390 29 397 31
rect 390 27 393 29
rect 395 27 397 29
rect 390 25 397 27
rect 405 30 412 32
rect 405 28 407 30
rect 409 28 412 30
rect 405 26 412 28
rect 414 26 423 39
rect 390 21 395 25
rect 416 22 423 26
rect 359 19 362 21
rect 364 19 366 21
rect 359 17 366 19
rect 379 19 381 21
rect 383 19 386 21
rect 379 17 386 19
rect 416 20 418 22
rect 420 20 423 22
rect 416 17 423 20
rect 425 30 433 39
rect 425 28 428 30
rect 430 28 433 30
rect 425 17 433 28
rect 435 37 443 39
rect 435 35 438 37
rect 440 35 443 37
rect 435 30 443 35
rect 435 28 438 30
rect 440 28 443 30
rect 435 23 443 28
rect 435 21 438 23
rect 440 21 443 23
rect 435 17 443 21
rect 445 37 457 39
rect 445 35 452 37
rect 454 35 457 37
rect 445 17 457 35
rect 459 29 464 39
rect 468 37 475 39
rect 468 35 470 37
rect 472 35 475 37
rect 468 33 475 35
rect 459 21 466 29
rect 470 26 475 33
rect 477 31 486 39
rect 507 32 512 39
rect 477 26 488 31
rect 479 21 488 26
rect 490 29 497 31
rect 490 27 493 29
rect 495 27 497 29
rect 490 25 497 27
rect 505 30 512 32
rect 505 28 507 30
rect 509 28 512 30
rect 505 26 512 28
rect 514 26 523 39
rect 490 21 495 25
rect 516 22 523 26
rect 459 19 462 21
rect 464 19 466 21
rect 459 17 466 19
rect 479 19 481 21
rect 483 19 486 21
rect 479 17 486 19
rect 516 20 518 22
rect 520 20 523 22
rect 516 17 523 20
rect 525 30 533 39
rect 525 28 528 30
rect 530 28 533 30
rect 525 17 533 28
rect 535 37 543 39
rect 535 35 538 37
rect 540 35 543 37
rect 535 30 543 35
rect 535 28 538 30
rect 540 28 543 30
rect 535 23 543 28
rect 535 21 538 23
rect 540 21 543 23
rect 535 17 543 21
rect 545 37 557 39
rect 545 35 552 37
rect 554 35 557 37
rect 545 17 557 35
rect 559 29 564 39
rect 568 37 575 39
rect 568 35 570 37
rect 572 35 575 37
rect 568 33 575 35
rect 559 21 566 29
rect 570 26 575 33
rect 577 31 586 39
rect 607 32 612 39
rect 577 26 588 31
rect 579 21 588 26
rect 590 29 597 31
rect 590 27 593 29
rect 595 27 597 29
rect 590 25 597 27
rect 605 30 612 32
rect 605 28 607 30
rect 609 28 612 30
rect 605 26 612 28
rect 614 26 623 39
rect 590 21 595 25
rect 616 22 623 26
rect 559 19 562 21
rect 564 19 566 21
rect 559 17 566 19
rect 579 19 581 21
rect 583 19 586 21
rect 579 17 586 19
rect 616 20 618 22
rect 620 20 623 22
rect 616 17 623 20
rect 625 30 633 39
rect 625 28 628 30
rect 630 28 633 30
rect 625 17 633 28
rect 635 37 643 39
rect 635 35 638 37
rect 640 35 643 37
rect 635 30 643 35
rect 635 28 638 30
rect 640 28 643 30
rect 635 23 643 28
rect 635 21 638 23
rect 640 21 643 23
rect 635 17 643 21
rect 645 37 657 39
rect 645 35 652 37
rect 654 35 657 37
rect 645 17 657 35
rect 659 29 664 39
rect 668 37 675 39
rect 668 35 670 37
rect 672 35 675 37
rect 668 33 675 35
rect 659 21 666 29
rect 670 26 675 33
rect 677 31 686 39
rect 707 32 712 39
rect 677 26 688 31
rect 679 21 688 26
rect 690 29 697 31
rect 690 27 693 29
rect 695 27 697 29
rect 690 25 697 27
rect 705 30 712 32
rect 705 28 707 30
rect 709 28 712 30
rect 705 26 712 28
rect 714 26 723 39
rect 690 21 695 25
rect 716 22 723 26
rect 659 19 662 21
rect 664 19 666 21
rect 659 17 666 19
rect 679 19 681 21
rect 683 19 686 21
rect 679 17 686 19
rect 716 20 718 22
rect 720 20 723 22
rect 716 17 723 20
rect 725 30 733 39
rect 725 28 728 30
rect 730 28 733 30
rect 725 17 733 28
rect 735 37 743 39
rect 735 35 738 37
rect 740 35 743 37
rect 735 30 743 35
rect 735 28 738 30
rect 740 28 743 30
rect 735 23 743 28
rect 735 21 738 23
rect 740 21 743 23
rect 735 17 743 21
rect 745 37 757 39
rect 745 35 752 37
rect 754 35 757 37
rect 745 17 757 35
rect 759 29 764 39
rect 768 37 775 39
rect 768 35 770 37
rect 772 35 775 37
rect 768 33 775 35
rect 759 21 766 29
rect 770 26 775 33
rect 777 31 786 39
rect 777 26 788 31
rect 779 21 788 26
rect 790 29 797 31
rect 790 27 793 29
rect 795 27 797 29
rect 790 25 797 27
rect 790 21 795 25
rect 759 19 762 21
rect 764 19 766 21
rect 759 17 766 19
rect 779 19 781 21
rect 783 19 786 21
rect 779 17 786 19
rect -1 -38 6 -35
rect -1 -40 1 -38
rect 3 -40 6 -38
rect -1 -44 6 -40
rect -12 -46 -5 -44
rect -12 -48 -10 -46
rect -8 -48 -5 -46
rect -12 -50 -5 -48
rect -10 -57 -5 -50
rect -3 -57 6 -44
rect 8 -46 16 -35
rect 8 -48 11 -46
rect 13 -48 16 -46
rect 8 -57 16 -48
rect 18 -39 26 -35
rect 18 -41 21 -39
rect 23 -41 26 -39
rect 18 -46 26 -41
rect 18 -48 21 -46
rect 23 -48 26 -46
rect 18 -53 26 -48
rect 18 -55 21 -53
rect 23 -55 26 -53
rect 18 -57 26 -55
rect 28 -53 40 -35
rect 28 -55 35 -53
rect 37 -55 40 -53
rect 28 -57 40 -55
rect 42 -37 49 -35
rect 42 -39 45 -37
rect 47 -39 49 -37
rect 62 -37 69 -35
rect 62 -39 64 -37
rect 66 -39 69 -37
rect 105 -38 112 -35
rect 42 -47 49 -39
rect 62 -44 71 -39
rect 42 -57 47 -47
rect 53 -51 58 -44
rect 51 -53 58 -51
rect 51 -55 53 -53
rect 55 -55 58 -53
rect 51 -57 58 -55
rect 60 -49 71 -44
rect 73 -43 78 -39
rect 73 -45 80 -43
rect 105 -40 107 -38
rect 109 -40 112 -38
rect 105 -44 112 -40
rect 73 -47 76 -45
rect 78 -47 80 -45
rect 73 -49 80 -47
rect 94 -46 101 -44
rect 94 -48 96 -46
rect 98 -48 101 -46
rect 60 -57 69 -49
rect 94 -50 101 -48
rect 96 -57 101 -50
rect 103 -57 112 -44
rect 114 -46 122 -35
rect 114 -48 117 -46
rect 119 -48 122 -46
rect 114 -57 122 -48
rect 124 -39 132 -35
rect 124 -41 127 -39
rect 129 -41 132 -39
rect 124 -46 132 -41
rect 124 -48 127 -46
rect 129 -48 132 -46
rect 124 -53 132 -48
rect 124 -55 127 -53
rect 129 -55 132 -53
rect 124 -57 132 -55
rect 134 -53 146 -35
rect 134 -55 141 -53
rect 143 -55 146 -53
rect 134 -57 146 -55
rect 148 -37 155 -35
rect 148 -39 151 -37
rect 153 -39 155 -37
rect 168 -37 175 -35
rect 168 -39 170 -37
rect 172 -39 175 -37
rect 211 -38 218 -35
rect 148 -47 155 -39
rect 168 -44 177 -39
rect 148 -57 153 -47
rect 159 -51 164 -44
rect 157 -53 164 -51
rect 157 -55 159 -53
rect 161 -55 164 -53
rect 157 -57 164 -55
rect 166 -49 177 -44
rect 179 -43 184 -39
rect 179 -45 186 -43
rect 211 -40 213 -38
rect 215 -40 218 -38
rect 211 -44 218 -40
rect 179 -47 182 -45
rect 184 -47 186 -45
rect 179 -49 186 -47
rect 200 -46 207 -44
rect 200 -48 202 -46
rect 204 -48 207 -46
rect 166 -57 175 -49
rect 200 -50 207 -48
rect 202 -57 207 -50
rect 209 -57 218 -44
rect 220 -46 228 -35
rect 220 -48 223 -46
rect 225 -48 228 -46
rect 220 -57 228 -48
rect 230 -39 238 -35
rect 230 -41 233 -39
rect 235 -41 238 -39
rect 230 -46 238 -41
rect 230 -48 233 -46
rect 235 -48 238 -46
rect 230 -53 238 -48
rect 230 -55 233 -53
rect 235 -55 238 -53
rect 230 -57 238 -55
rect 240 -53 252 -35
rect 240 -55 247 -53
rect 249 -55 252 -53
rect 240 -57 252 -55
rect 254 -37 261 -35
rect 254 -39 257 -37
rect 259 -39 261 -37
rect 274 -37 281 -35
rect 274 -39 276 -37
rect 278 -39 281 -37
rect 317 -38 324 -35
rect 254 -47 261 -39
rect 274 -44 283 -39
rect 254 -57 259 -47
rect 265 -51 270 -44
rect 263 -53 270 -51
rect 263 -55 265 -53
rect 267 -55 270 -53
rect 263 -57 270 -55
rect 272 -49 283 -44
rect 285 -43 290 -39
rect 285 -45 292 -43
rect 317 -40 319 -38
rect 321 -40 324 -38
rect 317 -44 324 -40
rect 285 -47 288 -45
rect 290 -47 292 -45
rect 285 -49 292 -47
rect 306 -46 313 -44
rect 306 -48 308 -46
rect 310 -48 313 -46
rect 272 -57 281 -49
rect 306 -50 313 -48
rect 308 -57 313 -50
rect 315 -57 324 -44
rect 326 -46 334 -35
rect 326 -48 329 -46
rect 331 -48 334 -46
rect 326 -57 334 -48
rect 336 -39 344 -35
rect 336 -41 339 -39
rect 341 -41 344 -39
rect 336 -46 344 -41
rect 336 -48 339 -46
rect 341 -48 344 -46
rect 336 -53 344 -48
rect 336 -55 339 -53
rect 341 -55 344 -53
rect 336 -57 344 -55
rect 346 -53 358 -35
rect 346 -55 353 -53
rect 355 -55 358 -53
rect 346 -57 358 -55
rect 360 -37 367 -35
rect 360 -39 363 -37
rect 365 -39 367 -37
rect 380 -37 387 -35
rect 380 -39 382 -37
rect 384 -39 387 -37
rect 423 -38 430 -35
rect 360 -47 367 -39
rect 380 -44 389 -39
rect 360 -57 365 -47
rect 371 -51 376 -44
rect 369 -53 376 -51
rect 369 -55 371 -53
rect 373 -55 376 -53
rect 369 -57 376 -55
rect 378 -49 389 -44
rect 391 -43 396 -39
rect 391 -45 398 -43
rect 423 -40 425 -38
rect 427 -40 430 -38
rect 423 -44 430 -40
rect 391 -47 394 -45
rect 396 -47 398 -45
rect 391 -49 398 -47
rect 412 -46 419 -44
rect 412 -48 414 -46
rect 416 -48 419 -46
rect 378 -57 387 -49
rect 412 -50 419 -48
rect 414 -57 419 -50
rect 421 -57 430 -44
rect 432 -46 440 -35
rect 432 -48 435 -46
rect 437 -48 440 -46
rect 432 -57 440 -48
rect 442 -39 450 -35
rect 442 -41 445 -39
rect 447 -41 450 -39
rect 442 -46 450 -41
rect 442 -48 445 -46
rect 447 -48 450 -46
rect 442 -53 450 -48
rect 442 -55 445 -53
rect 447 -55 450 -53
rect 442 -57 450 -55
rect 452 -53 464 -35
rect 452 -55 459 -53
rect 461 -55 464 -53
rect 452 -57 464 -55
rect 466 -37 473 -35
rect 466 -39 469 -37
rect 471 -39 473 -37
rect 486 -37 493 -35
rect 486 -39 488 -37
rect 490 -39 493 -37
rect 529 -38 536 -35
rect 466 -47 473 -39
rect 486 -44 495 -39
rect 466 -57 471 -47
rect 477 -51 482 -44
rect 475 -53 482 -51
rect 475 -55 477 -53
rect 479 -55 482 -53
rect 475 -57 482 -55
rect 484 -49 495 -44
rect 497 -43 502 -39
rect 497 -45 504 -43
rect 529 -40 531 -38
rect 533 -40 536 -38
rect 529 -44 536 -40
rect 497 -47 500 -45
rect 502 -47 504 -45
rect 497 -49 504 -47
rect 518 -46 525 -44
rect 518 -48 520 -46
rect 522 -48 525 -46
rect 484 -57 493 -49
rect 518 -50 525 -48
rect 520 -57 525 -50
rect 527 -57 536 -44
rect 538 -46 546 -35
rect 538 -48 541 -46
rect 543 -48 546 -46
rect 538 -57 546 -48
rect 548 -39 556 -35
rect 548 -41 551 -39
rect 553 -41 556 -39
rect 548 -46 556 -41
rect 548 -48 551 -46
rect 553 -48 556 -46
rect 548 -53 556 -48
rect 548 -55 551 -53
rect 553 -55 556 -53
rect 548 -57 556 -55
rect 558 -53 570 -35
rect 558 -55 565 -53
rect 567 -55 570 -53
rect 558 -57 570 -55
rect 572 -37 579 -35
rect 572 -39 575 -37
rect 577 -39 579 -37
rect 592 -37 599 -35
rect 592 -39 594 -37
rect 596 -39 599 -37
rect 635 -38 642 -35
rect 572 -47 579 -39
rect 592 -44 601 -39
rect 572 -57 577 -47
rect 583 -51 588 -44
rect 581 -53 588 -51
rect 581 -55 583 -53
rect 585 -55 588 -53
rect 581 -57 588 -55
rect 590 -49 601 -44
rect 603 -43 608 -39
rect 603 -45 610 -43
rect 635 -40 637 -38
rect 639 -40 642 -38
rect 635 -44 642 -40
rect 603 -47 606 -45
rect 608 -47 610 -45
rect 603 -49 610 -47
rect 624 -46 631 -44
rect 624 -48 626 -46
rect 628 -48 631 -46
rect 590 -57 599 -49
rect 624 -50 631 -48
rect 626 -57 631 -50
rect 633 -57 642 -44
rect 644 -46 652 -35
rect 644 -48 647 -46
rect 649 -48 652 -46
rect 644 -57 652 -48
rect 654 -39 662 -35
rect 654 -41 657 -39
rect 659 -41 662 -39
rect 654 -46 662 -41
rect 654 -48 657 -46
rect 659 -48 662 -46
rect 654 -53 662 -48
rect 654 -55 657 -53
rect 659 -55 662 -53
rect 654 -57 662 -55
rect 664 -53 676 -35
rect 664 -55 671 -53
rect 673 -55 676 -53
rect 664 -57 676 -55
rect 678 -37 685 -35
rect 678 -39 681 -37
rect 683 -39 685 -37
rect 698 -37 705 -35
rect 698 -39 700 -37
rect 702 -39 705 -37
rect 741 -38 748 -35
rect 678 -47 685 -39
rect 698 -44 707 -39
rect 678 -57 683 -47
rect 689 -51 694 -44
rect 687 -53 694 -51
rect 687 -55 689 -53
rect 691 -55 694 -53
rect 687 -57 694 -55
rect 696 -49 707 -44
rect 709 -43 714 -39
rect 709 -45 716 -43
rect 741 -40 743 -38
rect 745 -40 748 -38
rect 741 -44 748 -40
rect 709 -47 712 -45
rect 714 -47 716 -45
rect 709 -49 716 -47
rect 730 -46 737 -44
rect 730 -48 732 -46
rect 734 -48 737 -46
rect 696 -57 705 -49
rect 730 -50 737 -48
rect 732 -57 737 -50
rect 739 -57 748 -44
rect 750 -46 758 -35
rect 750 -48 753 -46
rect 755 -48 758 -46
rect 750 -57 758 -48
rect 760 -39 768 -35
rect 760 -41 763 -39
rect 765 -41 768 -39
rect 760 -46 768 -41
rect 760 -48 763 -46
rect 765 -48 768 -46
rect 760 -53 768 -48
rect 760 -55 763 -53
rect 765 -55 768 -53
rect 760 -57 768 -55
rect 770 -53 782 -35
rect 770 -55 777 -53
rect 779 -55 782 -53
rect 770 -57 782 -55
rect 784 -37 791 -35
rect 784 -39 787 -37
rect 789 -39 791 -37
rect 804 -37 811 -35
rect 804 -39 806 -37
rect 808 -39 811 -37
rect 847 -38 854 -35
rect 784 -47 791 -39
rect 804 -44 813 -39
rect 784 -57 789 -47
rect 795 -51 800 -44
rect 793 -53 800 -51
rect 793 -55 795 -53
rect 797 -55 800 -53
rect 793 -57 800 -55
rect 802 -49 813 -44
rect 815 -43 820 -39
rect 815 -45 822 -43
rect 847 -40 849 -38
rect 851 -40 854 -38
rect 847 -44 854 -40
rect 815 -47 818 -45
rect 820 -47 822 -45
rect 815 -49 822 -47
rect 836 -46 843 -44
rect 836 -48 838 -46
rect 840 -48 843 -46
rect 802 -57 811 -49
rect 836 -50 843 -48
rect 838 -57 843 -50
rect 845 -57 854 -44
rect 856 -46 864 -35
rect 856 -48 859 -46
rect 861 -48 864 -46
rect 856 -57 864 -48
rect 866 -39 874 -35
rect 866 -41 869 -39
rect 871 -41 874 -39
rect 866 -46 874 -41
rect 866 -48 869 -46
rect 871 -48 874 -46
rect 866 -53 874 -48
rect 866 -55 869 -53
rect 871 -55 874 -53
rect 866 -57 874 -55
rect 876 -53 888 -35
rect 876 -55 883 -53
rect 885 -55 888 -53
rect 876 -57 888 -55
rect 890 -37 897 -35
rect 890 -39 893 -37
rect 895 -39 897 -37
rect 910 -37 917 -35
rect 910 -39 912 -37
rect 914 -39 917 -37
rect 890 -47 897 -39
rect 910 -44 919 -39
rect 890 -57 895 -47
rect 901 -51 906 -44
rect 899 -53 906 -51
rect 899 -55 901 -53
rect 903 -55 906 -53
rect 899 -57 906 -55
rect 908 -49 919 -44
rect 921 -43 926 -39
rect 921 -45 928 -43
rect 921 -47 924 -45
rect 926 -47 928 -45
rect 921 -49 928 -47
rect 908 -57 917 -49
<< alu1 >>
rect 76 1183 385 1188
rect 76 1181 83 1183
rect 85 1181 136 1183
rect 138 1181 150 1183
rect 152 1181 171 1183
rect 173 1181 187 1183
rect 189 1181 197 1183
rect 199 1181 231 1183
rect 233 1181 284 1183
rect 286 1181 338 1183
rect 340 1181 361 1183
rect 363 1181 373 1183
rect 375 1181 385 1183
rect 76 1180 385 1181
rect 563 1183 747 1188
rect 563 1181 569 1183
rect 571 1181 589 1183
rect 591 1181 607 1183
rect 609 1181 660 1183
rect 662 1181 678 1183
rect 680 1181 690 1183
rect 692 1181 702 1183
rect 704 1181 747 1183
rect 563 1180 747 1181
rect 148 1174 165 1175
rect 116 1173 140 1174
rect 116 1171 118 1173
rect 120 1171 140 1173
rect 116 1170 140 1171
rect 88 1165 101 1167
rect 88 1163 89 1165
rect 91 1163 101 1165
rect 88 1162 101 1163
rect 136 1166 140 1170
rect 88 1161 98 1162
rect 96 1160 98 1161
rect 100 1160 101 1162
rect 80 1149 85 1151
rect 80 1147 82 1149
rect 84 1147 85 1149
rect 80 1142 85 1147
rect 96 1153 101 1160
rect 136 1164 137 1166
rect 139 1164 140 1166
rect 80 1140 81 1142
rect 83 1140 85 1142
rect 80 1135 85 1140
rect 80 1129 92 1135
rect 136 1142 140 1164
rect 124 1141 140 1142
rect 124 1140 133 1141
rect 124 1138 126 1140
rect 128 1139 133 1140
rect 135 1139 140 1141
rect 128 1138 140 1139
rect 124 1137 140 1138
rect 148 1172 161 1174
rect 163 1172 165 1174
rect 148 1171 165 1172
rect 148 1169 160 1171
rect 148 1141 152 1169
rect 184 1172 196 1175
rect 298 1174 310 1175
rect 184 1171 193 1172
rect 184 1169 186 1171
rect 188 1170 193 1171
rect 195 1170 196 1172
rect 188 1169 196 1170
rect 264 1173 288 1174
rect 164 1166 168 1167
rect 164 1164 165 1166
rect 167 1164 168 1166
rect 164 1161 168 1164
rect 164 1160 176 1161
rect 156 1157 160 1159
rect 164 1158 167 1160
rect 169 1158 176 1160
rect 164 1157 176 1158
rect 156 1155 157 1157
rect 159 1155 160 1157
rect 156 1153 160 1155
rect 172 1153 176 1157
rect 156 1149 168 1153
rect 164 1147 165 1149
rect 167 1147 168 1149
rect 164 1145 168 1147
rect 184 1149 188 1169
rect 264 1171 266 1173
rect 268 1171 288 1173
rect 264 1170 288 1171
rect 208 1163 213 1167
rect 208 1161 210 1163
rect 212 1161 213 1163
rect 208 1158 213 1161
rect 184 1147 189 1149
rect 184 1145 186 1147
rect 188 1145 189 1147
rect 148 1140 157 1141
rect 148 1138 153 1140
rect 155 1138 157 1140
rect 148 1137 157 1138
rect 151 1136 157 1137
rect 184 1140 189 1145
rect 184 1138 186 1140
rect 188 1138 189 1140
rect 199 1157 213 1158
rect 199 1155 203 1157
rect 205 1155 213 1157
rect 199 1154 213 1155
rect 236 1166 249 1167
rect 236 1164 237 1166
rect 239 1164 249 1166
rect 236 1162 249 1164
rect 236 1161 246 1162
rect 244 1160 246 1161
rect 248 1160 249 1162
rect 207 1149 220 1150
rect 207 1147 213 1149
rect 215 1147 220 1149
rect 207 1146 220 1147
rect 184 1136 189 1138
rect 151 1134 154 1136
rect 156 1134 157 1136
rect 151 1133 157 1134
rect 151 1131 153 1133
rect 155 1131 157 1133
rect 151 1130 157 1131
rect 216 1140 220 1146
rect 216 1138 217 1140
rect 219 1138 220 1140
rect 216 1137 220 1138
rect 228 1149 233 1151
rect 228 1147 230 1149
rect 232 1147 233 1149
rect 228 1135 233 1147
rect 244 1153 249 1160
rect 284 1163 288 1170
rect 284 1161 285 1163
rect 287 1161 288 1163
rect 228 1132 240 1135
rect 228 1130 235 1132
rect 237 1130 240 1132
rect 228 1129 240 1130
rect 284 1142 288 1161
rect 272 1140 288 1142
rect 272 1138 274 1140
rect 276 1138 288 1140
rect 272 1137 288 1138
rect 298 1172 299 1174
rect 301 1172 306 1174
rect 308 1172 310 1174
rect 298 1171 310 1172
rect 298 1143 302 1171
rect 314 1167 318 1175
rect 306 1163 318 1167
rect 322 1166 326 1175
rect 330 1169 342 1175
rect 322 1164 323 1166
rect 325 1164 326 1166
rect 306 1160 310 1163
rect 306 1158 307 1160
rect 309 1158 310 1160
rect 322 1159 326 1164
rect 338 1163 342 1169
rect 338 1161 339 1163
rect 341 1161 342 1163
rect 306 1157 310 1158
rect 306 1155 307 1157
rect 309 1155 310 1157
rect 306 1153 310 1155
rect 314 1155 326 1159
rect 314 1150 320 1155
rect 314 1148 317 1150
rect 319 1148 320 1150
rect 314 1145 320 1148
rect 330 1149 334 1159
rect 338 1157 342 1161
rect 338 1155 339 1157
rect 341 1155 342 1157
rect 338 1153 342 1155
rect 358 1166 362 1175
rect 640 1173 664 1174
rect 358 1164 360 1166
rect 330 1148 342 1149
rect 330 1146 339 1148
rect 341 1146 342 1148
rect 330 1145 342 1146
rect 298 1141 310 1143
rect 298 1140 334 1141
rect 298 1138 310 1140
rect 312 1138 330 1140
rect 332 1138 334 1140
rect 298 1137 334 1138
rect 329 1133 334 1137
rect 329 1131 330 1133
rect 332 1131 334 1133
rect 329 1129 334 1131
rect 338 1129 342 1145
rect 358 1148 362 1164
rect 640 1171 642 1173
rect 644 1171 664 1173
rect 640 1170 664 1171
rect 366 1159 370 1167
rect 566 1166 586 1167
rect 566 1164 579 1166
rect 581 1164 586 1166
rect 566 1161 586 1164
rect 366 1158 378 1159
rect 366 1157 374 1158
rect 366 1155 367 1157
rect 369 1156 374 1157
rect 376 1156 378 1158
rect 369 1155 378 1156
rect 366 1153 378 1155
rect 358 1146 360 1148
rect 358 1143 362 1146
rect 358 1141 370 1143
rect 358 1139 360 1141
rect 362 1140 370 1141
rect 362 1139 367 1140
rect 358 1138 367 1139
rect 369 1138 370 1140
rect 566 1142 570 1161
rect 590 1156 594 1159
rect 592 1154 594 1156
rect 612 1162 625 1167
rect 612 1161 622 1162
rect 620 1160 622 1161
rect 624 1160 625 1162
rect 590 1150 594 1154
rect 581 1149 594 1150
rect 581 1147 591 1149
rect 593 1147 594 1149
rect 581 1146 594 1147
rect 604 1149 609 1151
rect 604 1147 606 1149
rect 608 1147 609 1149
rect 566 1141 583 1142
rect 566 1139 574 1141
rect 576 1139 579 1141
rect 581 1139 583 1141
rect 566 1138 583 1139
rect 358 1137 370 1138
rect 604 1135 609 1147
rect 620 1156 625 1160
rect 660 1162 664 1170
rect 660 1160 661 1162
rect 663 1160 664 1162
rect 620 1154 621 1156
rect 623 1154 625 1156
rect 620 1153 625 1154
rect 604 1132 616 1135
rect 604 1130 605 1132
rect 607 1130 616 1132
rect 604 1129 616 1130
rect 660 1142 664 1160
rect 648 1140 664 1142
rect 648 1138 650 1140
rect 652 1138 664 1140
rect 648 1137 664 1138
rect 675 1166 679 1175
rect 675 1164 677 1166
rect 675 1148 679 1164
rect 683 1166 687 1167
rect 683 1164 684 1166
rect 686 1164 687 1166
rect 706 1166 711 1175
rect 725 1173 743 1174
rect 725 1171 727 1173
rect 729 1171 730 1173
rect 732 1171 743 1173
rect 725 1170 743 1171
rect 706 1165 733 1166
rect 683 1159 687 1164
rect 706 1163 708 1165
rect 710 1163 730 1165
rect 732 1163 733 1165
rect 706 1162 733 1163
rect 729 1160 730 1162
rect 732 1160 733 1162
rect 683 1157 695 1159
rect 729 1158 733 1160
rect 683 1155 684 1157
rect 686 1155 695 1157
rect 683 1153 695 1155
rect 706 1157 723 1158
rect 706 1155 719 1157
rect 721 1155 723 1157
rect 706 1154 723 1155
rect 675 1146 677 1148
rect 675 1143 679 1146
rect 706 1148 711 1154
rect 739 1150 743 1170
rect 706 1146 707 1148
rect 709 1146 711 1148
rect 706 1145 711 1146
rect 721 1149 743 1150
rect 721 1147 740 1149
rect 742 1147 743 1149
rect 721 1145 722 1147
rect 724 1146 743 1147
rect 724 1145 727 1146
rect 675 1142 687 1143
rect 675 1141 682 1142
rect 675 1139 677 1141
rect 679 1140 682 1141
rect 684 1140 687 1142
rect 679 1139 687 1140
rect 675 1137 687 1139
rect 721 1140 727 1145
rect 721 1138 722 1140
rect 724 1138 727 1140
rect 721 1136 727 1138
rect 76 1123 385 1124
rect 76 1121 116 1123
rect 118 1121 187 1123
rect 189 1121 264 1123
rect 266 1121 341 1123
rect 343 1121 361 1123
rect 363 1121 373 1123
rect 375 1121 385 1123
rect 76 1116 385 1121
rect 563 1123 747 1124
rect 563 1121 588 1123
rect 590 1121 640 1123
rect 642 1121 678 1123
rect 680 1121 690 1123
rect 692 1121 747 1123
rect 76 1111 336 1116
rect 76 1109 119 1111
rect 121 1109 131 1111
rect 133 1109 147 1111
rect 149 1109 221 1111
rect 223 1109 235 1111
rect 237 1109 261 1111
rect 263 1109 301 1111
rect 303 1109 323 1111
rect 325 1109 336 1111
rect 76 1108 336 1109
rect 563 1111 747 1121
rect 563 1109 572 1111
rect 574 1109 584 1111
rect 586 1109 604 1111
rect 606 1109 705 1111
rect 707 1109 747 1111
rect 563 1108 747 1109
rect 80 1089 92 1095
rect 116 1093 128 1095
rect 116 1091 118 1093
rect 120 1091 128 1093
rect 116 1089 128 1091
rect 144 1094 149 1096
rect 144 1092 146 1094
rect 148 1092 149 1094
rect 188 1095 193 1103
rect 144 1091 149 1092
rect 144 1089 145 1091
rect 147 1089 149 1091
rect 80 1070 84 1089
rect 96 1086 108 1087
rect 96 1084 105 1086
rect 107 1084 108 1086
rect 96 1081 108 1084
rect 80 1068 81 1070
rect 83 1068 84 1070
rect 80 1061 84 1068
rect 88 1077 92 1079
rect 106 1079 108 1081
rect 88 1075 89 1077
rect 91 1075 92 1077
rect 88 1071 92 1075
rect 104 1073 108 1079
rect 116 1086 120 1089
rect 116 1084 118 1086
rect 88 1068 100 1071
rect 88 1066 97 1068
rect 99 1066 100 1068
rect 88 1065 100 1066
rect 116 1068 120 1084
rect 144 1087 149 1089
rect 144 1085 146 1087
rect 148 1085 149 1087
rect 144 1083 149 1085
rect 124 1078 136 1079
rect 124 1077 133 1078
rect 124 1075 125 1077
rect 127 1076 133 1077
rect 135 1076 136 1078
rect 127 1075 136 1076
rect 124 1073 136 1075
rect 116 1066 118 1068
rect 80 1060 89 1061
rect 80 1058 85 1060
rect 87 1058 89 1060
rect 80 1057 89 1058
rect 116 1060 120 1066
rect 124 1065 128 1073
rect 116 1058 117 1060
rect 119 1058 120 1060
rect 116 1057 120 1058
rect 144 1063 148 1083
rect 176 1086 180 1095
rect 167 1085 180 1086
rect 167 1083 168 1085
rect 170 1083 173 1085
rect 175 1083 180 1085
rect 167 1082 180 1083
rect 188 1093 190 1095
rect 192 1094 193 1095
rect 192 1093 201 1094
rect 188 1091 198 1093
rect 200 1091 201 1093
rect 188 1090 201 1091
rect 188 1088 192 1090
rect 188 1086 190 1088
rect 159 1077 173 1078
rect 159 1075 163 1077
rect 165 1075 173 1077
rect 159 1074 173 1075
rect 168 1071 173 1074
rect 144 1061 146 1063
rect 148 1061 156 1063
rect 144 1057 156 1061
rect 168 1069 169 1071
rect 171 1069 173 1071
rect 168 1065 173 1069
rect 188 1067 192 1086
rect 219 1086 225 1094
rect 256 1101 316 1102
rect 256 1099 257 1101
rect 259 1099 316 1101
rect 256 1098 316 1099
rect 211 1085 233 1086
rect 211 1084 221 1085
rect 211 1082 217 1084
rect 219 1083 221 1084
rect 223 1083 233 1085
rect 219 1082 233 1083
rect 256 1078 260 1098
rect 264 1093 297 1094
rect 264 1091 265 1093
rect 267 1091 293 1093
rect 295 1091 297 1093
rect 264 1090 297 1091
rect 203 1077 216 1078
rect 203 1075 207 1077
rect 209 1075 216 1077
rect 203 1074 216 1075
rect 188 1065 190 1067
rect 188 1057 192 1065
rect 212 1068 216 1074
rect 227 1077 233 1078
rect 227 1075 229 1077
rect 231 1075 233 1077
rect 227 1071 233 1075
rect 256 1076 258 1078
rect 256 1074 260 1076
rect 212 1066 213 1068
rect 215 1066 216 1068
rect 212 1065 216 1066
rect 220 1068 233 1071
rect 220 1066 230 1068
rect 232 1066 233 1068
rect 220 1065 233 1066
rect 264 1062 268 1090
rect 312 1086 316 1098
rect 577 1093 589 1095
rect 577 1091 582 1093
rect 584 1091 585 1093
rect 587 1091 589 1093
rect 577 1089 589 1091
rect 272 1085 307 1086
rect 272 1083 273 1085
rect 275 1083 307 1085
rect 272 1082 307 1083
rect 312 1082 327 1086
rect 585 1086 589 1089
rect 587 1084 589 1086
rect 272 1071 276 1082
rect 303 1078 307 1082
rect 321 1078 327 1082
rect 272 1069 273 1071
rect 275 1069 276 1071
rect 287 1070 293 1078
rect 303 1074 316 1078
rect 321 1076 323 1078
rect 325 1076 327 1078
rect 321 1075 327 1076
rect 569 1077 581 1079
rect 569 1076 578 1077
rect 312 1072 316 1074
rect 569 1074 574 1076
rect 576 1075 578 1076
rect 580 1075 581 1077
rect 576 1074 581 1075
rect 569 1073 581 1074
rect 312 1070 313 1072
rect 315 1070 316 1072
rect 272 1067 276 1069
rect 282 1069 307 1070
rect 282 1067 284 1069
rect 286 1067 298 1069
rect 300 1067 303 1069
rect 305 1067 307 1069
rect 312 1068 316 1070
rect 320 1070 324 1071
rect 320 1068 321 1070
rect 323 1068 324 1070
rect 282 1066 307 1067
rect 320 1063 324 1068
rect 264 1060 294 1062
rect 264 1058 268 1060
rect 270 1058 290 1060
rect 292 1058 294 1060
rect 264 1057 294 1058
rect 312 1061 324 1063
rect 312 1059 313 1061
rect 315 1059 324 1061
rect 312 1057 324 1059
rect 577 1065 581 1073
rect 585 1068 589 1084
rect 587 1066 589 1068
rect 585 1057 589 1066
rect 601 1094 606 1096
rect 601 1092 603 1094
rect 605 1092 606 1094
rect 601 1087 606 1092
rect 601 1085 603 1087
rect 605 1085 606 1087
rect 601 1083 606 1085
rect 633 1094 637 1095
rect 633 1092 634 1094
rect 636 1092 637 1094
rect 601 1081 602 1083
rect 604 1081 605 1083
rect 601 1063 605 1081
rect 633 1086 637 1092
rect 663 1089 675 1095
rect 624 1085 637 1086
rect 624 1083 630 1085
rect 632 1083 637 1085
rect 624 1082 637 1083
rect 647 1086 659 1087
rect 647 1084 655 1086
rect 657 1084 659 1086
rect 647 1081 659 1084
rect 647 1079 649 1081
rect 616 1077 630 1078
rect 616 1075 620 1077
rect 622 1075 630 1077
rect 616 1074 630 1075
rect 601 1061 603 1063
rect 605 1061 613 1063
rect 601 1057 613 1061
rect 625 1068 630 1074
rect 647 1073 651 1079
rect 663 1077 667 1079
rect 663 1075 664 1077
rect 666 1075 667 1077
rect 663 1071 667 1075
rect 625 1066 627 1068
rect 629 1066 630 1068
rect 625 1065 630 1066
rect 655 1069 667 1071
rect 655 1067 664 1069
rect 666 1067 667 1069
rect 655 1065 667 1067
rect 671 1061 675 1089
rect 666 1060 675 1061
rect 666 1058 668 1060
rect 670 1058 672 1060
rect 674 1058 675 1060
rect 683 1094 699 1095
rect 683 1092 691 1094
rect 693 1092 695 1094
rect 697 1092 699 1094
rect 683 1090 699 1092
rect 683 1069 687 1090
rect 731 1097 743 1103
rect 738 1093 743 1097
rect 738 1091 740 1093
rect 742 1091 743 1093
rect 683 1067 684 1069
rect 686 1067 687 1069
rect 683 1062 687 1067
rect 722 1072 727 1079
rect 738 1085 743 1091
rect 738 1083 739 1085
rect 741 1083 743 1085
rect 738 1081 743 1083
rect 722 1070 723 1072
rect 725 1071 727 1072
rect 725 1070 735 1071
rect 722 1068 735 1070
rect 722 1066 732 1068
rect 734 1066 735 1068
rect 722 1065 735 1066
rect 683 1061 707 1062
rect 683 1059 703 1061
rect 705 1059 707 1061
rect 683 1058 707 1059
rect 666 1057 675 1058
rect 76 1051 336 1052
rect 76 1049 119 1051
rect 121 1049 131 1051
rect 133 1049 147 1051
rect 149 1049 157 1051
rect 159 1049 191 1051
rect 193 1049 201 1051
rect 203 1049 279 1051
rect 281 1049 323 1051
rect 325 1049 336 1051
rect 76 1044 336 1049
rect 563 1051 747 1052
rect 563 1049 572 1051
rect 574 1049 584 1051
rect 586 1049 604 1051
rect 606 1049 614 1051
rect 616 1049 685 1051
rect 687 1049 738 1051
rect 740 1049 747 1051
rect 563 1044 747 1049
rect 76 1039 308 1044
rect 76 1037 83 1039
rect 85 1037 136 1039
rect 138 1037 195 1039
rect 197 1037 211 1039
rect 213 1037 233 1039
rect 235 1037 293 1039
rect 295 1037 303 1039
rect 305 1037 308 1039
rect 76 1036 308 1037
rect 507 1039 747 1044
rect 507 1037 514 1039
rect 516 1037 526 1039
rect 528 1037 578 1039
rect 580 1037 648 1039
rect 650 1037 658 1039
rect 660 1037 676 1039
rect 678 1037 688 1039
rect 690 1037 702 1039
rect 704 1037 747 1039
rect 507 1036 747 1037
rect 148 1030 157 1031
rect 116 1029 140 1030
rect 116 1027 118 1029
rect 120 1027 140 1029
rect 116 1026 140 1027
rect 88 1021 101 1023
rect 88 1019 89 1021
rect 91 1019 101 1021
rect 88 1018 101 1019
rect 88 1017 98 1018
rect 96 1016 98 1017
rect 100 1016 101 1018
rect 80 1005 85 1007
rect 80 1003 82 1005
rect 84 1003 85 1005
rect 80 998 85 1003
rect 96 1009 101 1016
rect 136 1020 140 1026
rect 136 1018 137 1020
rect 139 1018 140 1020
rect 80 996 81 998
rect 83 996 85 998
rect 80 991 85 996
rect 80 985 92 991
rect 136 998 140 1018
rect 124 996 140 998
rect 124 994 126 996
rect 128 994 140 996
rect 124 993 140 994
rect 148 1028 153 1030
rect 155 1028 157 1030
rect 148 1027 157 1028
rect 148 999 152 1027
rect 203 1029 216 1031
rect 203 1027 204 1029
rect 206 1027 216 1029
rect 220 1030 248 1031
rect 220 1028 222 1030
rect 224 1028 244 1030
rect 246 1028 248 1030
rect 220 1027 248 1028
rect 203 1026 216 1027
rect 156 1020 168 1023
rect 211 1022 216 1026
rect 156 1018 161 1020
rect 163 1018 168 1020
rect 195 1021 207 1022
rect 195 1019 196 1021
rect 198 1019 207 1021
rect 195 1018 204 1019
rect 156 1017 168 1018
rect 203 1017 204 1018
rect 206 1017 207 1019
rect 211 1021 219 1022
rect 211 1019 215 1021
rect 217 1019 219 1021
rect 211 1018 219 1019
rect 226 1021 232 1023
rect 226 1019 227 1021
rect 229 1019 232 1021
rect 156 1013 160 1017
rect 156 1011 157 1013
rect 159 1011 160 1013
rect 156 1009 160 1011
rect 172 1009 176 1015
rect 203 1014 207 1017
rect 226 1014 232 1019
rect 192 1013 199 1014
rect 192 1011 194 1013
rect 196 1011 199 1013
rect 192 1010 199 1011
rect 203 1010 232 1014
rect 236 1021 240 1023
rect 236 1019 237 1021
rect 239 1019 240 1021
rect 174 1007 176 1009
rect 164 1004 176 1007
rect 164 1002 168 1004
rect 170 1002 176 1004
rect 195 1006 199 1010
rect 236 1006 240 1019
rect 195 1005 240 1006
rect 195 1003 237 1005
rect 239 1003 240 1005
rect 195 1002 240 1003
rect 164 1001 176 1002
rect 148 996 160 999
rect 244 998 248 1027
rect 304 1029 308 1031
rect 304 1027 305 1029
rect 307 1027 308 1029
rect 263 1021 276 1023
rect 263 1019 273 1021
rect 275 1019 276 1021
rect 263 1017 276 1019
rect 263 1013 269 1017
rect 263 1011 265 1013
rect 267 1011 269 1013
rect 263 1010 269 1011
rect 280 1014 284 1023
rect 304 1023 308 1027
rect 306 1021 308 1023
rect 280 1013 293 1014
rect 280 1011 287 1013
rect 289 1011 290 1013
rect 292 1011 293 1013
rect 280 1010 293 1011
rect 263 1004 277 1006
rect 279 1004 285 1006
rect 263 1002 285 1004
rect 148 994 149 996
rect 151 994 160 996
rect 211 997 248 998
rect 211 996 245 997
rect 211 994 218 996
rect 220 995 245 996
rect 247 995 248 997
rect 220 994 248 995
rect 148 993 160 994
rect 271 997 277 1002
rect 271 995 272 997
rect 274 995 277 997
rect 271 994 277 995
rect 304 1002 308 1021
rect 306 1000 308 1002
rect 304 998 308 1000
rect 295 995 308 998
rect 295 994 304 995
rect 303 993 304 994
rect 306 993 308 995
rect 511 1030 515 1031
rect 511 1028 512 1030
rect 514 1028 515 1030
rect 511 1022 515 1028
rect 511 1020 513 1022
rect 511 1004 515 1020
rect 519 1015 523 1023
rect 582 1022 587 1031
rect 601 1029 619 1030
rect 601 1027 603 1029
rect 605 1027 619 1029
rect 601 1026 619 1027
rect 582 1021 609 1022
rect 582 1019 584 1021
rect 586 1019 606 1021
rect 608 1019 609 1021
rect 582 1018 609 1019
rect 605 1016 606 1018
rect 608 1016 609 1018
rect 519 1014 531 1015
rect 605 1014 609 1016
rect 519 1013 528 1014
rect 519 1011 520 1013
rect 522 1012 528 1013
rect 530 1012 531 1014
rect 522 1011 531 1012
rect 519 1009 531 1011
rect 555 1013 599 1014
rect 555 1011 556 1013
rect 558 1011 595 1013
rect 597 1011 599 1013
rect 555 1010 599 1011
rect 511 1002 513 1004
rect 511 999 515 1002
rect 582 1001 587 1010
rect 615 1006 619 1026
rect 634 1021 639 1023
rect 634 1019 636 1021
rect 638 1019 639 1021
rect 634 1014 639 1019
rect 651 1027 663 1031
rect 651 1025 659 1027
rect 661 1025 663 1027
rect 634 1013 648 1014
rect 634 1011 642 1013
rect 644 1011 648 1013
rect 634 1010 648 1011
rect 597 1003 619 1006
rect 597 1001 598 1003
rect 600 1002 619 1003
rect 627 1005 640 1006
rect 627 1003 628 1005
rect 630 1003 632 1005
rect 634 1003 640 1005
rect 627 1002 640 1003
rect 600 1001 603 1002
rect 597 999 603 1001
rect 511 997 523 999
rect 511 995 513 997
rect 515 995 523 997
rect 511 993 523 995
rect 597 997 598 999
rect 600 997 603 999
rect 597 996 603 997
rect 597 994 598 996
rect 600 994 603 996
rect 303 985 308 993
rect 597 992 603 994
rect 627 993 631 1002
rect 659 1005 663 1025
rect 658 1003 663 1005
rect 658 1001 659 1003
rect 661 1001 663 1003
rect 658 998 663 1001
rect 673 1022 677 1031
rect 673 1020 675 1022
rect 673 1004 677 1020
rect 681 1015 685 1023
rect 706 1022 711 1031
rect 725 1029 743 1030
rect 725 1027 727 1029
rect 729 1027 743 1029
rect 725 1026 743 1027
rect 706 1021 733 1022
rect 706 1019 708 1021
rect 710 1019 715 1021
rect 717 1019 733 1021
rect 706 1018 733 1019
rect 729 1016 730 1018
rect 732 1016 733 1018
rect 681 1013 693 1015
rect 729 1014 733 1016
rect 681 1011 682 1013
rect 684 1011 688 1013
rect 690 1011 693 1013
rect 681 1009 693 1011
rect 706 1013 723 1014
rect 706 1011 719 1013
rect 721 1011 723 1013
rect 706 1010 723 1011
rect 673 1002 675 1004
rect 673 1001 677 1002
rect 673 999 674 1001
rect 676 999 677 1001
rect 706 1004 711 1010
rect 739 1006 743 1026
rect 706 1002 707 1004
rect 709 1002 711 1004
rect 706 1001 711 1002
rect 721 1003 743 1006
rect 721 1001 722 1003
rect 724 1002 743 1003
rect 724 1001 727 1002
rect 721 1000 727 1001
rect 658 997 666 998
rect 658 996 663 997
rect 658 994 659 996
rect 661 995 663 996
rect 665 995 666 997
rect 661 994 666 995
rect 673 997 685 999
rect 673 995 675 997
rect 677 995 685 997
rect 658 992 663 994
rect 673 993 685 995
rect 721 998 724 1000
rect 726 998 727 1000
rect 721 996 727 998
rect 721 994 722 996
rect 724 994 727 996
rect 721 992 727 994
rect 76 979 308 980
rect 76 977 116 979
rect 118 977 259 979
rect 261 977 273 979
rect 275 977 308 979
rect 76 967 308 977
rect 76 965 119 967
rect 121 965 131 967
rect 133 965 147 967
rect 149 965 222 967
rect 224 965 299 967
rect 301 965 308 967
rect 76 964 308 965
rect 507 979 747 980
rect 507 977 514 979
rect 516 977 526 979
rect 528 977 658 979
rect 660 977 676 979
rect 678 977 688 979
rect 690 977 747 979
rect 507 967 747 977
rect 507 965 533 967
rect 535 965 582 967
rect 584 965 626 967
rect 628 965 634 967
rect 636 965 705 967
rect 707 965 747 967
rect 507 964 747 965
rect 83 957 89 958
rect 83 955 85 957
rect 87 955 89 957
rect 83 951 89 955
rect 80 950 89 951
rect 80 948 85 950
rect 87 948 89 950
rect 80 947 89 948
rect 116 949 128 951
rect 116 947 118 949
rect 120 947 128 949
rect 80 924 84 947
rect 116 945 128 947
rect 144 950 149 952
rect 144 948 146 950
rect 148 948 149 950
rect 96 942 108 943
rect 96 940 105 942
rect 107 940 108 942
rect 96 939 108 940
rect 116 942 120 945
rect 116 940 118 942
rect 88 935 100 939
rect 88 933 92 935
rect 88 931 89 933
rect 91 931 92 933
rect 104 934 108 935
rect 104 932 105 934
rect 107 932 108 934
rect 104 931 108 932
rect 88 929 92 931
rect 96 930 108 931
rect 80 922 81 924
rect 83 922 84 924
rect 80 919 84 922
rect 96 928 99 930
rect 101 928 108 930
rect 96 927 108 928
rect 96 921 100 927
rect 116 924 120 940
rect 144 943 149 948
rect 144 941 146 943
rect 148 941 149 943
rect 144 939 149 941
rect 176 949 180 951
rect 176 947 177 949
rect 179 947 180 949
rect 124 933 136 935
rect 124 931 125 933
rect 127 931 136 933
rect 124 929 136 931
rect 116 922 118 924
rect 80 917 92 919
rect 77 916 99 917
rect 77 914 78 916
rect 80 914 93 916
rect 95 914 99 916
rect 77 913 99 914
rect 116 916 120 922
rect 124 924 128 929
rect 124 922 125 924
rect 127 922 128 924
rect 144 925 148 939
rect 144 923 145 925
rect 147 923 148 925
rect 124 921 128 922
rect 116 914 117 916
rect 119 914 120 916
rect 116 913 120 914
rect 144 919 148 923
rect 176 942 180 947
rect 167 941 180 942
rect 167 939 173 941
rect 175 939 180 941
rect 167 938 180 939
rect 200 950 216 951
rect 200 948 212 950
rect 214 948 216 950
rect 200 946 216 948
rect 200 934 204 946
rect 248 957 260 959
rect 248 955 249 957
rect 251 955 260 957
rect 248 953 260 955
rect 159 933 173 934
rect 159 931 163 933
rect 165 931 173 933
rect 159 930 173 931
rect 168 926 173 930
rect 200 932 201 934
rect 203 932 204 934
rect 144 917 146 919
rect 148 917 156 919
rect 144 913 156 917
rect 168 921 189 926
rect 184 916 189 921
rect 184 914 185 916
rect 187 914 189 916
rect 200 918 204 932
rect 239 928 244 935
rect 255 941 260 953
rect 255 939 256 941
rect 258 939 260 941
rect 255 937 260 939
rect 268 950 272 951
rect 268 948 269 950
rect 271 948 272 950
rect 268 942 272 948
rect 299 950 304 952
rect 268 941 281 942
rect 268 939 273 941
rect 275 939 281 941
rect 268 938 281 939
rect 239 926 240 928
rect 242 927 244 928
rect 242 926 252 927
rect 239 925 252 926
rect 239 923 240 925
rect 242 923 252 925
rect 239 921 252 923
rect 275 933 289 934
rect 275 931 283 933
rect 285 931 289 933
rect 275 930 289 931
rect 299 948 300 950
rect 302 948 304 950
rect 299 946 304 948
rect 299 944 300 946
rect 302 944 304 946
rect 299 943 304 944
rect 299 941 300 943
rect 302 941 304 943
rect 299 939 304 941
rect 275 924 280 930
rect 275 922 277 924
rect 279 922 280 924
rect 275 921 280 922
rect 200 917 224 918
rect 200 915 220 917
rect 222 915 224 917
rect 300 919 304 939
rect 200 914 224 915
rect 292 917 300 919
rect 302 917 304 919
rect 184 913 189 914
rect 292 913 304 917
rect 511 950 527 951
rect 511 948 523 950
rect 525 948 527 950
rect 511 946 527 948
rect 511 926 515 946
rect 559 958 571 959
rect 559 956 567 958
rect 569 956 571 958
rect 559 953 571 956
rect 511 924 512 926
rect 514 924 515 926
rect 511 918 515 924
rect 550 928 555 935
rect 566 941 571 953
rect 566 939 567 941
rect 569 939 571 941
rect 566 937 571 939
rect 579 950 584 952
rect 579 948 581 950
rect 583 948 584 950
rect 579 943 584 948
rect 579 941 581 943
rect 583 941 584 943
rect 579 939 584 941
rect 611 949 615 951
rect 611 947 612 949
rect 614 947 615 949
rect 550 926 551 928
rect 553 927 555 928
rect 553 926 563 927
rect 550 925 563 926
rect 550 923 558 925
rect 560 923 563 925
rect 550 921 563 923
rect 579 925 583 939
rect 579 923 580 925
rect 582 923 583 925
rect 511 917 535 918
rect 511 915 531 917
rect 533 915 535 917
rect 579 919 583 923
rect 611 942 615 947
rect 635 950 639 952
rect 635 948 636 950
rect 638 948 639 950
rect 635 943 639 948
rect 655 950 659 952
rect 655 948 656 950
rect 658 948 659 950
rect 602 941 615 942
rect 602 939 608 941
rect 610 939 615 941
rect 602 938 615 939
rect 623 934 627 943
rect 635 941 636 943
rect 638 942 639 943
rect 655 943 659 948
rect 683 950 699 951
rect 683 949 695 950
rect 683 947 689 949
rect 691 948 695 949
rect 697 948 699 950
rect 691 947 699 948
rect 683 946 699 947
rect 655 942 656 943
rect 638 941 656 942
rect 658 941 659 943
rect 635 939 644 941
rect 646 939 659 941
rect 635 938 659 939
rect 594 933 608 934
rect 594 931 598 933
rect 600 931 605 933
rect 607 931 608 933
rect 594 930 608 931
rect 579 917 581 919
rect 583 917 591 919
rect 511 914 535 915
rect 579 913 591 917
rect 603 921 608 930
rect 623 933 636 934
rect 623 931 627 933
rect 629 931 632 933
rect 634 931 636 933
rect 623 929 636 931
rect 655 924 659 938
rect 663 934 675 935
rect 663 933 672 934
rect 663 931 664 933
rect 666 932 672 933
rect 674 932 675 934
rect 666 931 675 932
rect 663 929 675 931
rect 655 922 656 924
rect 658 922 659 924
rect 655 920 659 922
rect 671 921 675 929
rect 683 918 687 946
rect 731 953 743 959
rect 738 949 743 953
rect 738 947 740 949
rect 742 947 743 949
rect 722 928 727 935
rect 738 941 743 947
rect 738 939 739 941
rect 741 939 743 941
rect 738 937 743 939
rect 722 926 723 928
rect 725 927 727 928
rect 725 926 735 927
rect 722 925 735 926
rect 722 923 732 925
rect 734 923 735 925
rect 722 921 735 923
rect 683 917 707 918
rect 683 915 684 917
rect 686 915 703 917
rect 705 915 707 917
rect 683 914 707 915
rect 76 907 308 908
rect 76 905 82 907
rect 84 905 103 907
rect 105 905 119 907
rect 121 905 131 907
rect 133 905 147 907
rect 149 905 157 907
rect 159 905 202 907
rect 204 905 255 907
rect 257 905 289 907
rect 291 905 299 907
rect 301 905 308 907
rect 76 900 308 905
rect 507 907 747 908
rect 507 905 513 907
rect 515 905 566 907
rect 568 905 582 907
rect 584 905 592 907
rect 594 905 626 907
rect 628 905 685 907
rect 687 905 738 907
rect 740 905 747 907
rect 507 900 747 905
rect 76 895 392 900
rect 76 893 119 895
rect 121 893 129 895
rect 131 893 168 895
rect 170 893 178 895
rect 180 893 239 895
rect 241 893 249 895
rect 251 893 267 895
rect 269 893 279 895
rect 281 893 295 895
rect 297 893 305 895
rect 307 893 339 895
rect 341 893 349 895
rect 351 893 392 895
rect 76 892 392 893
rect 483 895 747 900
rect 483 893 507 895
rect 509 893 517 895
rect 519 893 534 895
rect 536 893 546 895
rect 548 893 580 895
rect 582 893 590 895
rect 592 893 610 895
rect 612 893 620 895
rect 622 893 684 895
rect 686 893 694 895
rect 696 893 747 895
rect 483 892 711 893
rect 713 892 747 893
rect 89 879 93 887
rect 104 885 109 887
rect 104 883 105 885
rect 107 883 109 885
rect 104 881 109 883
rect 77 878 93 879
rect 77 876 78 878
rect 80 876 93 878
rect 77 874 87 876
rect 89 874 93 876
rect 77 873 93 874
rect 105 878 109 881
rect 105 876 106 878
rect 108 876 109 878
rect 97 869 101 871
rect 97 867 98 869
rect 100 867 101 869
rect 97 866 101 867
rect 88 865 101 866
rect 88 863 97 865
rect 99 863 101 865
rect 88 862 101 863
rect 88 858 94 862
rect 105 854 109 876
rect 96 850 109 854
rect 116 883 128 887
rect 116 881 118 883
rect 120 881 128 883
rect 165 883 177 887
rect 116 861 120 881
rect 165 881 167 883
rect 169 881 177 883
rect 140 878 145 879
rect 140 876 141 878
rect 143 876 145 878
rect 140 870 145 876
rect 116 859 121 861
rect 116 857 118 859
rect 120 857 121 859
rect 116 852 121 857
rect 116 850 118 852
rect 120 850 121 852
rect 131 869 145 870
rect 131 867 135 869
rect 137 867 145 869
rect 131 866 145 867
rect 139 861 152 862
rect 139 859 140 861
rect 142 859 145 861
rect 147 859 152 861
rect 139 858 152 859
rect 116 847 121 850
rect 116 845 117 847
rect 119 845 121 847
rect 116 844 121 845
rect 148 849 152 858
rect 165 861 169 881
rect 189 875 194 879
rect 189 873 190 875
rect 192 873 194 875
rect 189 870 194 873
rect 165 859 170 861
rect 165 857 167 859
rect 169 857 170 859
rect 165 856 170 857
rect 165 854 166 856
rect 168 854 170 856
rect 165 852 170 854
rect 165 850 167 852
rect 169 850 170 852
rect 180 869 194 870
rect 180 867 184 869
rect 186 867 194 869
rect 180 866 194 867
rect 225 870 230 879
rect 242 883 254 887
rect 242 881 250 883
rect 252 881 254 883
rect 225 869 239 870
rect 225 867 229 869
rect 231 867 233 869
rect 235 867 239 869
rect 225 866 239 867
rect 188 861 201 862
rect 188 859 194 861
rect 196 859 201 861
rect 188 858 201 859
rect 165 848 170 850
rect 197 852 201 858
rect 197 850 198 852
rect 200 850 201 852
rect 197 849 201 850
rect 218 861 231 862
rect 218 859 223 861
rect 225 859 231 861
rect 218 858 231 859
rect 218 853 222 858
rect 250 864 254 881
rect 250 862 251 864
rect 253 862 254 864
rect 250 861 254 862
rect 218 851 219 853
rect 221 851 222 853
rect 218 849 222 851
rect 249 859 254 861
rect 249 857 250 859
rect 252 857 254 859
rect 249 852 254 857
rect 249 850 250 852
rect 252 850 254 852
rect 249 848 254 850
rect 264 878 268 887
rect 264 876 266 878
rect 264 875 268 876
rect 264 873 265 875
rect 267 873 268 875
rect 264 860 268 873
rect 272 871 276 879
rect 292 883 304 887
rect 292 881 294 883
rect 296 881 304 883
rect 272 869 284 871
rect 272 867 273 869
rect 275 868 284 869
rect 275 867 281 868
rect 272 866 281 867
rect 283 866 284 868
rect 272 865 284 866
rect 264 858 266 860
rect 264 855 268 858
rect 292 861 296 881
rect 336 879 340 887
rect 316 878 321 879
rect 316 876 317 878
rect 319 876 321 878
rect 316 870 321 876
rect 292 859 297 861
rect 292 857 294 859
rect 296 857 297 859
rect 292 856 297 857
rect 264 853 276 855
rect 264 851 266 853
rect 268 851 276 853
rect 264 849 276 851
rect 292 854 293 856
rect 295 854 297 856
rect 292 852 297 854
rect 292 850 294 852
rect 296 850 297 852
rect 307 869 321 870
rect 307 867 311 869
rect 313 867 321 869
rect 307 866 321 867
rect 336 877 338 879
rect 315 861 328 862
rect 315 859 321 861
rect 323 859 325 861
rect 327 859 328 861
rect 315 858 328 859
rect 292 848 297 850
rect 324 849 328 858
rect 336 858 340 877
rect 360 870 364 879
rect 368 878 381 879
rect 368 876 378 878
rect 380 876 381 878
rect 368 873 381 876
rect 351 869 364 870
rect 351 867 355 869
rect 357 867 361 869
rect 363 867 364 869
rect 351 866 364 867
rect 375 869 381 873
rect 375 867 377 869
rect 379 867 381 869
rect 375 866 381 867
rect 493 870 498 879
rect 510 883 522 887
rect 510 881 518 883
rect 520 881 522 883
rect 518 878 522 881
rect 493 869 507 870
rect 493 867 501 869
rect 503 867 504 869
rect 506 867 507 869
rect 493 866 507 867
rect 336 856 338 858
rect 336 854 340 856
rect 359 860 365 862
rect 367 860 381 862
rect 359 858 381 860
rect 486 861 499 862
rect 486 859 491 861
rect 493 859 499 861
rect 486 858 499 859
rect 336 851 349 854
rect 336 849 338 851
rect 340 850 349 851
rect 340 849 341 850
rect 336 845 341 849
rect 336 843 338 845
rect 340 843 341 845
rect 336 841 341 843
rect 367 853 373 858
rect 367 851 370 853
rect 372 851 373 853
rect 367 850 373 851
rect 486 852 490 858
rect 518 876 519 878
rect 521 876 522 878
rect 518 861 522 876
rect 486 850 487 852
rect 489 850 490 852
rect 486 849 490 850
rect 517 859 522 861
rect 517 857 518 859
rect 520 857 522 859
rect 517 852 522 857
rect 517 850 518 852
rect 520 850 522 852
rect 517 848 522 850
rect 531 878 535 887
rect 531 876 533 878
rect 531 860 535 876
rect 539 878 543 879
rect 539 876 540 878
rect 542 876 543 878
rect 566 878 571 879
rect 539 871 543 876
rect 566 876 567 878
rect 569 876 571 878
rect 539 869 551 871
rect 539 867 540 869
rect 542 867 551 869
rect 539 865 551 867
rect 566 870 571 876
rect 583 883 595 887
rect 583 881 591 883
rect 593 881 595 883
rect 566 869 580 870
rect 566 867 574 869
rect 576 867 580 869
rect 566 866 580 867
rect 531 858 533 860
rect 531 855 535 858
rect 559 861 572 862
rect 559 860 564 861
rect 559 858 560 860
rect 562 859 564 860
rect 566 859 572 861
rect 562 858 572 859
rect 531 853 543 855
rect 531 851 533 853
rect 535 852 543 853
rect 535 851 540 852
rect 531 850 540 851
rect 542 850 543 852
rect 531 849 543 850
rect 559 849 563 858
rect 591 861 595 881
rect 590 859 595 861
rect 590 857 591 859
rect 593 857 595 859
rect 590 855 595 857
rect 590 853 592 855
rect 594 853 595 855
rect 590 852 595 853
rect 590 850 591 852
rect 593 850 595 852
rect 590 848 595 850
rect 607 883 619 887
rect 607 881 609 883
rect 611 881 619 883
rect 607 861 611 881
rect 631 870 636 879
rect 607 859 612 861
rect 607 857 609 859
rect 611 857 612 859
rect 607 855 612 857
rect 607 853 609 855
rect 611 853 612 855
rect 607 852 612 853
rect 607 850 609 852
rect 611 850 612 852
rect 622 869 636 870
rect 622 867 623 869
rect 625 867 626 869
rect 628 867 636 869
rect 622 866 636 867
rect 654 873 667 879
rect 654 871 655 873
rect 657 871 660 873
rect 654 869 660 871
rect 654 867 656 869
rect 658 867 660 869
rect 654 866 660 867
rect 671 870 675 879
rect 695 879 699 887
rect 703 886 711 887
rect 703 884 704 886
rect 706 884 711 886
rect 703 883 711 884
rect 734 886 743 887
rect 734 884 736 886
rect 738 884 743 886
rect 734 883 743 884
rect 697 877 699 879
rect 671 869 684 870
rect 671 867 678 869
rect 680 867 681 869
rect 683 867 684 869
rect 671 866 684 867
rect 630 861 643 862
rect 630 859 636 861
rect 638 859 643 861
rect 630 858 643 859
rect 654 860 668 862
rect 670 860 676 862
rect 654 858 676 860
rect 695 867 699 877
rect 695 865 696 867
rect 698 865 699 867
rect 707 870 711 883
rect 722 877 735 879
rect 722 875 724 877
rect 726 875 735 877
rect 722 874 735 875
rect 707 869 720 870
rect 707 867 712 869
rect 714 867 720 869
rect 707 866 720 867
rect 731 869 735 874
rect 731 867 732 869
rect 734 867 735 869
rect 731 865 735 867
rect 607 848 612 850
rect 639 852 643 858
rect 639 850 640 852
rect 642 850 643 852
rect 639 849 643 850
rect 662 854 668 858
rect 662 852 664 854
rect 666 852 668 854
rect 662 850 668 852
rect 695 858 699 865
rect 697 856 699 858
rect 695 854 699 856
rect 686 851 699 854
rect 686 850 695 851
rect 694 849 695 850
rect 697 849 699 851
rect 707 861 726 862
rect 707 859 722 861
rect 724 859 726 861
rect 707 858 726 859
rect 707 852 711 858
rect 739 854 743 883
rect 707 850 708 852
rect 710 850 711 852
rect 707 849 711 850
rect 718 852 743 854
rect 718 850 719 852
rect 721 850 739 852
rect 741 850 743 852
rect 718 849 722 850
rect 694 841 699 849
rect 718 847 719 849
rect 721 847 722 849
rect 718 845 722 847
rect 718 843 719 845
rect 721 843 722 845
rect 718 841 722 843
rect 738 845 743 850
rect 738 843 739 845
rect 741 843 743 845
rect 738 841 743 843
rect 76 835 392 836
rect 76 833 84 835
rect 86 833 92 835
rect 94 833 119 835
rect 121 833 168 835
rect 170 833 249 835
rect 251 833 267 835
rect 269 833 279 835
rect 281 833 295 835
rect 297 833 369 835
rect 371 833 383 835
rect 385 833 392 835
rect 76 828 392 833
rect 483 835 747 836
rect 483 833 517 835
rect 519 833 534 835
rect 536 833 546 835
rect 548 833 590 835
rect 592 833 610 835
rect 612 833 650 835
rect 652 833 664 835
rect 666 833 747 835
rect 483 828 747 833
rect 76 823 340 828
rect 76 821 157 823
rect 159 821 171 823
rect 173 821 211 823
rect 213 821 231 823
rect 233 821 275 823
rect 277 821 287 823
rect 289 821 304 823
rect 306 821 340 823
rect 76 820 340 821
rect 431 823 747 828
rect 431 821 438 823
rect 440 821 452 823
rect 454 821 526 823
rect 528 821 542 823
rect 544 821 554 823
rect 556 821 572 823
rect 574 821 653 823
rect 655 821 702 823
rect 704 821 729 823
rect 731 821 737 823
rect 739 821 747 823
rect 431 820 747 821
rect 80 813 85 815
rect 80 811 82 813
rect 84 811 85 813
rect 80 806 85 811
rect 101 813 105 815
rect 101 811 102 813
rect 104 811 105 813
rect 101 809 105 811
rect 101 807 102 809
rect 104 807 105 809
rect 124 807 129 815
rect 101 806 105 807
rect 80 804 82 806
rect 84 804 102 806
rect 104 804 105 806
rect 80 802 105 804
rect 112 806 116 807
rect 112 804 113 806
rect 115 804 116 806
rect 80 773 84 802
rect 112 798 116 804
rect 97 797 116 798
rect 97 795 99 797
rect 101 795 116 797
rect 97 794 116 795
rect 124 805 126 807
rect 128 806 129 807
rect 128 805 137 806
rect 124 802 137 805
rect 124 800 128 802
rect 124 798 126 800
rect 88 789 92 791
rect 88 787 89 789
rect 91 787 92 789
rect 88 782 92 787
rect 103 789 116 790
rect 103 787 109 789
rect 111 787 116 789
rect 103 786 116 787
rect 88 781 101 782
rect 88 779 97 781
rect 99 779 101 781
rect 88 777 101 779
rect 112 773 116 786
rect 124 779 128 798
rect 155 804 161 806
rect 155 802 157 804
rect 159 802 161 804
rect 155 798 161 802
rect 180 806 184 807
rect 180 804 181 806
rect 183 804 184 806
rect 180 798 184 804
rect 211 806 216 808
rect 147 796 169 798
rect 147 794 153 796
rect 155 794 169 796
rect 180 797 193 798
rect 180 795 185 797
rect 187 795 193 797
rect 180 794 193 795
rect 139 789 152 790
rect 139 787 140 789
rect 142 787 143 789
rect 145 787 152 789
rect 139 786 152 787
rect 124 777 126 779
rect 80 772 89 773
rect 80 770 85 772
rect 87 770 89 772
rect 80 769 89 770
rect 112 772 120 773
rect 112 770 117 772
rect 119 770 120 772
rect 112 769 120 770
rect 124 772 128 777
rect 148 777 152 786
rect 163 789 169 790
rect 163 787 165 789
rect 167 787 169 789
rect 163 785 169 787
rect 163 783 166 785
rect 168 783 169 785
rect 156 777 169 783
rect 187 789 201 790
rect 187 787 195 789
rect 197 787 198 789
rect 200 787 201 789
rect 187 786 201 787
rect 211 804 212 806
rect 214 804 216 806
rect 211 803 216 804
rect 211 801 212 803
rect 214 801 216 803
rect 211 799 216 801
rect 211 797 212 799
rect 214 797 216 799
rect 211 795 216 797
rect 187 777 192 786
rect 124 770 125 772
rect 127 770 128 772
rect 124 769 128 770
rect 212 775 216 795
rect 204 773 212 775
rect 214 773 216 775
rect 204 769 216 773
rect 228 806 233 808
rect 228 804 230 806
rect 232 804 233 806
rect 228 803 233 804
rect 228 801 229 803
rect 231 801 233 803
rect 228 799 233 801
rect 228 797 230 799
rect 232 797 233 799
rect 228 795 233 797
rect 228 775 232 795
rect 260 798 264 807
rect 280 806 292 807
rect 280 804 281 806
rect 283 805 292 806
rect 283 804 288 805
rect 280 803 288 804
rect 290 803 292 805
rect 280 801 292 803
rect 251 797 261 798
rect 251 795 257 797
rect 259 796 261 797
rect 263 796 264 798
rect 259 795 264 796
rect 251 794 264 795
rect 288 798 292 801
rect 290 796 292 798
rect 243 789 257 790
rect 243 787 247 789
rect 249 787 257 789
rect 243 786 257 787
rect 228 773 230 775
rect 232 773 240 775
rect 228 769 240 773
rect 252 780 257 786
rect 272 789 284 791
rect 272 787 281 789
rect 283 787 284 789
rect 272 785 284 787
rect 252 778 254 780
rect 256 778 257 780
rect 280 780 284 785
rect 252 777 257 778
rect 280 778 281 780
rect 283 778 284 780
rect 280 777 284 778
rect 288 780 292 796
rect 290 778 292 780
rect 288 769 292 778
rect 301 806 306 808
rect 301 804 303 806
rect 305 804 306 806
rect 301 799 306 804
rect 301 797 303 799
rect 305 797 306 799
rect 301 795 306 797
rect 333 806 337 807
rect 333 804 334 806
rect 336 804 337 806
rect 301 780 305 795
rect 301 778 302 780
rect 304 778 305 780
rect 333 798 337 804
rect 450 805 456 806
rect 450 803 451 805
rect 453 803 456 805
rect 450 798 456 803
rect 482 813 487 815
rect 482 811 483 813
rect 485 811 487 813
rect 482 807 487 811
rect 482 806 483 807
rect 474 805 483 806
rect 485 805 487 807
rect 474 802 487 805
rect 324 797 337 798
rect 324 795 330 797
rect 332 795 337 797
rect 324 794 337 795
rect 442 796 464 798
rect 442 794 456 796
rect 458 794 464 796
rect 483 800 487 802
rect 485 798 487 800
rect 316 789 330 790
rect 316 787 317 789
rect 319 787 320 789
rect 322 787 330 789
rect 316 786 330 787
rect 301 775 305 778
rect 301 773 303 775
rect 305 773 313 775
rect 301 769 313 773
rect 325 777 330 786
rect 442 789 448 790
rect 442 787 444 789
rect 446 787 448 789
rect 442 783 448 787
rect 459 789 472 790
rect 459 787 460 789
rect 462 787 466 789
rect 468 787 472 789
rect 459 786 472 787
rect 442 780 455 783
rect 442 778 443 780
rect 445 778 455 780
rect 442 777 455 778
rect 459 777 463 786
rect 483 779 487 798
rect 495 798 499 807
rect 526 806 531 808
rect 495 797 508 798
rect 495 795 496 797
rect 498 795 500 797
rect 502 795 508 797
rect 495 794 508 795
rect 485 777 487 779
rect 502 789 516 790
rect 502 787 510 789
rect 512 787 516 789
rect 502 786 516 787
rect 526 804 527 806
rect 529 804 531 806
rect 526 802 531 804
rect 526 800 528 802
rect 530 800 531 802
rect 547 805 559 807
rect 547 803 555 805
rect 557 803 559 805
rect 547 801 559 803
rect 526 799 531 800
rect 526 797 527 799
rect 529 797 531 799
rect 526 795 531 797
rect 502 780 507 786
rect 502 778 504 780
rect 506 778 507 780
rect 502 777 507 778
rect 483 769 487 777
rect 527 775 531 795
rect 555 798 559 801
rect 557 796 559 798
rect 539 790 551 791
rect 539 788 540 790
rect 542 789 551 790
rect 542 788 548 789
rect 539 787 548 788
rect 550 787 551 789
rect 539 785 551 787
rect 519 773 527 775
rect 529 773 531 775
rect 519 769 531 773
rect 547 777 551 785
rect 555 783 559 796
rect 555 781 556 783
rect 558 781 559 783
rect 555 780 559 781
rect 557 778 559 780
rect 555 769 559 778
rect 569 806 574 808
rect 569 804 571 806
rect 573 804 574 806
rect 569 799 574 804
rect 569 797 571 799
rect 573 797 574 799
rect 569 795 574 797
rect 601 805 605 807
rect 601 803 602 805
rect 604 803 605 805
rect 569 794 573 795
rect 569 792 570 794
rect 572 792 573 794
rect 569 775 573 792
rect 601 798 605 803
rect 592 797 605 798
rect 592 795 598 797
rect 600 795 605 797
rect 592 794 605 795
rect 622 806 626 807
rect 622 804 623 806
rect 625 804 626 806
rect 622 798 626 804
rect 653 806 658 808
rect 622 797 635 798
rect 622 795 627 797
rect 629 795 635 797
rect 622 794 635 795
rect 584 789 598 790
rect 584 787 588 789
rect 590 787 592 789
rect 594 787 598 789
rect 584 786 598 787
rect 569 773 571 775
rect 573 773 581 775
rect 569 769 581 773
rect 593 777 598 786
rect 629 789 643 790
rect 629 787 637 789
rect 639 787 643 789
rect 629 786 643 787
rect 653 804 654 806
rect 656 804 658 806
rect 653 802 658 804
rect 653 800 655 802
rect 657 800 658 802
rect 653 799 658 800
rect 653 797 654 799
rect 656 797 658 799
rect 653 795 658 797
rect 629 783 634 786
rect 629 781 631 783
rect 633 781 634 783
rect 629 777 634 781
rect 654 775 658 795
rect 671 798 675 807
rect 702 811 707 812
rect 702 809 704 811
rect 706 809 707 811
rect 702 806 707 809
rect 671 797 684 798
rect 671 795 676 797
rect 678 795 681 797
rect 683 795 684 797
rect 671 794 684 795
rect 678 789 692 790
rect 678 787 686 789
rect 688 787 692 789
rect 678 786 692 787
rect 702 804 703 806
rect 705 804 707 806
rect 702 799 707 804
rect 702 797 703 799
rect 705 797 707 799
rect 702 795 707 797
rect 678 780 683 786
rect 678 778 680 780
rect 682 778 683 780
rect 678 777 683 778
rect 646 773 654 775
rect 656 773 658 775
rect 703 775 707 795
rect 646 769 658 773
rect 695 773 703 775
rect 705 773 707 775
rect 695 769 707 773
rect 714 802 727 806
rect 714 780 718 802
rect 729 794 735 798
rect 722 793 735 794
rect 722 791 724 793
rect 726 791 735 793
rect 722 790 735 791
rect 722 789 726 790
rect 722 787 723 789
rect 725 787 726 789
rect 722 785 726 787
rect 714 778 715 780
rect 717 778 718 780
rect 714 775 718 778
rect 730 782 746 783
rect 730 780 734 782
rect 736 780 746 782
rect 730 778 743 780
rect 745 778 746 780
rect 730 777 746 778
rect 714 773 719 775
rect 714 771 716 773
rect 718 771 719 773
rect 714 769 719 771
rect 730 769 734 777
rect 76 763 110 764
rect 112 763 340 764
rect 76 761 127 763
rect 129 761 137 763
rect 139 761 201 763
rect 203 761 211 763
rect 213 761 231 763
rect 233 761 241 763
rect 243 761 275 763
rect 277 761 287 763
rect 289 761 304 763
rect 306 761 314 763
rect 316 761 340 763
rect 76 756 340 761
rect 431 763 747 764
rect 431 761 472 763
rect 474 761 482 763
rect 484 761 516 763
rect 518 761 526 763
rect 528 761 542 763
rect 544 761 554 763
rect 556 761 572 763
rect 574 761 582 763
rect 584 761 643 763
rect 645 761 653 763
rect 655 761 692 763
rect 694 761 702 763
rect 704 761 747 763
rect 431 756 747 761
rect 76 751 344 756
rect 76 749 83 751
rect 85 749 136 751
rect 138 749 195 751
rect 197 749 229 751
rect 231 749 239 751
rect 241 749 255 751
rect 257 749 308 751
rect 310 749 323 751
rect 325 749 335 751
rect 337 749 344 751
rect 76 748 344 749
rect 515 751 747 756
rect 515 749 522 751
rect 524 749 532 751
rect 534 749 566 751
rect 568 749 619 751
rect 621 749 664 751
rect 666 749 674 751
rect 676 749 690 751
rect 692 749 702 751
rect 704 749 718 751
rect 720 749 739 751
rect 741 749 747 751
rect 515 748 747 749
rect 116 741 140 742
rect 116 739 118 741
rect 120 739 137 741
rect 139 739 140 741
rect 116 738 140 739
rect 88 733 101 735
rect 88 731 89 733
rect 91 731 101 733
rect 88 730 101 731
rect 88 729 98 730
rect 96 728 98 729
rect 100 728 101 730
rect 80 717 85 719
rect 80 715 82 717
rect 84 715 85 717
rect 80 711 85 715
rect 96 721 101 728
rect 80 709 81 711
rect 83 709 85 711
rect 80 703 85 709
rect 80 697 92 703
rect 136 710 140 738
rect 148 727 152 735
rect 164 734 168 736
rect 164 732 165 734
rect 167 732 168 734
rect 148 725 160 727
rect 148 724 157 725
rect 148 722 149 724
rect 151 723 157 724
rect 159 723 160 725
rect 151 722 160 723
rect 148 721 160 722
rect 164 718 168 732
rect 187 725 200 727
rect 187 723 189 725
rect 191 723 194 725
rect 196 723 200 725
rect 187 722 200 723
rect 215 726 220 735
rect 232 739 244 743
rect 288 741 312 742
rect 232 737 240 739
rect 242 737 244 739
rect 215 725 229 726
rect 215 723 216 725
rect 218 723 223 725
rect 225 723 229 725
rect 215 722 229 723
rect 164 717 188 718
rect 164 715 177 717
rect 179 715 188 717
rect 164 713 165 715
rect 167 714 185 715
rect 167 713 168 714
rect 124 709 140 710
rect 124 708 132 709
rect 124 706 126 708
rect 128 707 132 708
rect 134 707 140 709
rect 128 706 140 707
rect 124 705 140 706
rect 164 708 168 713
rect 184 713 185 714
rect 187 713 188 715
rect 196 713 200 722
rect 208 717 221 718
rect 208 715 213 717
rect 215 715 221 717
rect 208 714 221 715
rect 164 706 165 708
rect 167 706 168 708
rect 164 704 168 706
rect 184 708 188 713
rect 184 706 185 708
rect 187 706 188 708
rect 184 704 188 706
rect 208 709 212 714
rect 240 733 244 737
rect 288 739 290 741
rect 292 739 312 741
rect 288 738 312 739
rect 240 731 241 733
rect 243 731 244 733
rect 240 717 244 731
rect 260 733 273 735
rect 260 731 263 733
rect 265 731 273 733
rect 260 730 273 731
rect 260 729 270 730
rect 268 728 270 729
rect 272 728 273 730
rect 208 707 209 709
rect 211 707 212 709
rect 208 705 212 707
rect 239 715 244 717
rect 239 713 240 715
rect 242 713 244 715
rect 239 708 244 713
rect 239 706 240 708
rect 242 706 244 708
rect 239 704 244 706
rect 252 717 257 719
rect 252 715 254 717
rect 256 715 257 717
rect 252 703 257 715
rect 268 721 273 728
rect 308 731 312 738
rect 308 729 309 731
rect 311 729 312 731
rect 252 700 264 703
rect 252 698 254 700
rect 256 698 264 700
rect 252 697 264 698
rect 308 710 312 729
rect 296 708 312 710
rect 296 706 298 708
rect 300 706 312 708
rect 296 705 312 706
rect 320 734 324 743
rect 320 732 322 734
rect 320 716 324 732
rect 328 733 332 735
rect 519 739 531 743
rect 634 742 639 743
rect 519 737 521 739
rect 523 737 531 739
rect 599 741 623 742
rect 328 731 329 733
rect 331 731 332 733
rect 328 727 332 731
rect 328 725 340 727
rect 328 723 329 725
rect 331 723 340 725
rect 328 721 340 723
rect 320 714 322 716
rect 320 711 324 714
rect 519 717 523 737
rect 599 739 601 741
rect 603 739 623 741
rect 599 738 623 739
rect 543 734 548 735
rect 543 732 544 734
rect 546 732 548 734
rect 543 726 548 732
rect 519 715 524 717
rect 519 713 521 715
rect 523 713 524 715
rect 519 712 524 713
rect 320 709 332 711
rect 320 707 322 709
rect 324 707 329 709
rect 331 707 332 709
rect 320 705 332 707
rect 519 710 521 712
rect 523 710 524 712
rect 519 708 524 710
rect 519 706 521 708
rect 523 706 524 708
rect 534 725 548 726
rect 534 723 538 725
rect 540 723 548 725
rect 534 722 548 723
rect 571 733 584 735
rect 571 731 581 733
rect 583 731 584 733
rect 571 730 584 731
rect 571 729 581 730
rect 579 728 581 729
rect 583 728 584 730
rect 542 717 555 718
rect 542 715 548 717
rect 550 715 555 717
rect 542 714 555 715
rect 519 704 524 706
rect 551 708 555 714
rect 551 706 552 708
rect 554 706 555 708
rect 551 705 555 706
rect 563 717 568 719
rect 563 715 565 717
rect 567 715 568 717
rect 563 703 568 715
rect 579 721 584 728
rect 619 723 623 738
rect 634 740 636 742
rect 638 740 639 742
rect 634 735 639 740
rect 634 730 655 735
rect 667 739 679 743
rect 667 737 675 739
rect 677 737 679 739
rect 619 721 620 723
rect 622 721 623 723
rect 650 726 655 730
rect 650 725 664 726
rect 650 723 658 725
rect 660 723 664 725
rect 650 722 664 723
rect 563 701 575 703
rect 563 699 572 701
rect 574 699 575 701
rect 563 697 575 699
rect 619 710 623 721
rect 607 708 623 710
rect 607 706 609 708
rect 611 706 623 708
rect 607 705 623 706
rect 643 717 656 718
rect 643 715 648 717
rect 650 715 656 717
rect 643 714 656 715
rect 643 709 647 714
rect 675 733 679 737
rect 703 742 707 743
rect 703 740 704 742
rect 706 740 707 742
rect 695 734 699 735
rect 675 731 676 733
rect 678 731 679 733
rect 675 717 679 731
rect 695 732 696 734
rect 698 732 699 734
rect 695 727 699 732
rect 703 734 707 740
rect 724 742 746 743
rect 724 740 728 742
rect 730 740 743 742
rect 745 740 746 742
rect 724 739 746 740
rect 731 737 743 739
rect 705 732 707 734
rect 687 725 699 727
rect 687 723 696 725
rect 698 723 699 725
rect 687 721 699 723
rect 643 707 644 709
rect 646 707 647 709
rect 643 705 647 707
rect 674 715 679 717
rect 674 713 675 715
rect 677 713 679 715
rect 674 708 679 713
rect 703 716 707 732
rect 723 729 727 735
rect 715 728 727 729
rect 715 726 722 728
rect 724 726 727 728
rect 739 734 743 737
rect 739 732 740 734
rect 742 732 743 734
rect 715 725 727 726
rect 731 725 735 727
rect 715 724 719 725
rect 715 722 716 724
rect 718 722 719 724
rect 715 721 719 722
rect 731 723 732 725
rect 734 723 735 725
rect 731 721 735 723
rect 723 717 735 721
rect 705 714 707 716
rect 703 711 707 714
rect 715 716 727 717
rect 715 714 716 716
rect 718 714 727 716
rect 715 713 727 714
rect 674 706 675 708
rect 677 706 679 708
rect 674 704 679 706
rect 695 709 707 711
rect 739 709 743 732
rect 695 707 703 709
rect 705 707 707 709
rect 695 705 707 707
rect 734 708 743 709
rect 734 706 736 708
rect 738 706 743 708
rect 734 705 743 706
rect 734 701 740 705
rect 734 699 736 701
rect 738 699 740 701
rect 734 698 740 699
rect 76 691 344 692
rect 76 689 116 691
rect 118 689 187 691
rect 189 689 195 691
rect 197 689 239 691
rect 241 689 288 691
rect 290 689 323 691
rect 325 689 335 691
rect 337 689 344 691
rect 76 684 344 689
rect 515 691 747 692
rect 515 689 522 691
rect 524 689 599 691
rect 601 689 674 691
rect 676 689 690 691
rect 692 689 702 691
rect 704 689 747 691
rect 76 679 252 684
rect 76 677 133 679
rect 135 677 145 679
rect 147 677 163 679
rect 165 677 252 679
rect 76 676 252 677
rect 515 679 747 689
rect 515 677 548 679
rect 550 677 562 679
rect 564 677 705 679
rect 707 677 747 679
rect 515 676 747 677
rect 96 662 102 664
rect 96 660 99 662
rect 101 660 102 662
rect 96 658 102 660
rect 96 656 97 658
rect 99 656 102 658
rect 138 661 150 663
rect 160 662 165 664
rect 138 659 146 661
rect 148 659 150 661
rect 138 657 150 659
rect 157 661 162 662
rect 157 659 158 661
rect 160 660 162 661
rect 164 660 165 662
rect 160 659 165 660
rect 157 658 165 659
rect 96 655 102 656
rect 96 654 99 655
rect 80 653 99 654
rect 101 653 102 655
rect 80 650 102 653
rect 112 654 117 655
rect 112 652 114 654
rect 116 652 117 654
rect 80 630 84 650
rect 112 646 117 652
rect 146 655 147 657
rect 149 655 150 657
rect 146 654 150 655
rect 148 652 150 654
rect 100 645 117 646
rect 100 643 102 645
rect 104 643 117 645
rect 100 642 117 643
rect 130 645 142 647
rect 130 643 133 645
rect 135 643 139 645
rect 141 643 142 645
rect 90 640 94 642
rect 130 641 142 643
rect 90 638 91 640
rect 93 638 94 640
rect 90 637 117 638
rect 90 635 106 637
rect 108 635 113 637
rect 115 635 117 637
rect 90 634 117 635
rect 80 629 98 630
rect 80 627 94 629
rect 96 627 98 629
rect 80 626 98 627
rect 112 625 117 634
rect 138 633 142 641
rect 146 636 150 652
rect 148 634 150 636
rect 146 625 150 634
rect 160 655 165 658
rect 160 653 162 655
rect 164 653 165 655
rect 160 651 165 653
rect 160 631 164 651
rect 192 654 196 663
rect 220 662 226 664
rect 220 660 223 662
rect 225 660 226 662
rect 220 659 226 660
rect 220 657 223 659
rect 225 657 226 659
rect 220 655 226 657
rect 515 663 520 671
rect 515 661 517 663
rect 519 662 520 663
rect 519 661 528 662
rect 515 658 528 661
rect 515 656 519 658
rect 220 654 223 655
rect 183 653 196 654
rect 183 651 189 653
rect 191 651 193 653
rect 195 651 196 653
rect 183 650 196 651
rect 204 653 223 654
rect 225 653 226 655
rect 204 650 226 653
rect 175 645 189 646
rect 175 643 179 645
rect 181 643 189 645
rect 175 642 189 643
rect 160 629 162 631
rect 164 629 172 631
rect 160 625 172 629
rect 184 637 189 642
rect 184 635 185 637
rect 187 635 189 637
rect 184 633 189 635
rect 204 630 208 650
rect 236 646 241 655
rect 515 654 517 656
rect 224 645 268 646
rect 224 643 226 645
rect 228 643 265 645
rect 267 643 268 645
rect 224 642 268 643
rect 214 640 218 642
rect 214 638 215 640
rect 217 638 218 640
rect 214 637 241 638
rect 214 635 215 637
rect 217 635 237 637
rect 239 635 241 637
rect 214 634 241 635
rect 204 629 222 630
rect 204 627 218 629
rect 220 627 222 629
rect 204 626 222 627
rect 236 625 241 634
rect 515 635 519 654
rect 546 661 552 662
rect 546 659 549 661
rect 551 659 552 661
rect 546 654 552 659
rect 663 662 675 663
rect 575 661 603 662
rect 575 659 576 661
rect 578 660 603 661
rect 605 660 612 662
rect 578 659 612 660
rect 575 658 612 659
rect 663 660 672 662
rect 674 660 675 662
rect 538 652 560 654
rect 538 650 544 652
rect 546 650 560 652
rect 530 645 543 646
rect 530 643 531 645
rect 533 643 534 645
rect 536 643 543 645
rect 530 642 543 643
rect 515 633 517 635
rect 515 629 519 633
rect 539 633 543 642
rect 554 645 560 646
rect 554 643 556 645
rect 558 643 560 645
rect 554 639 560 643
rect 547 637 560 639
rect 547 635 548 637
rect 550 635 560 637
rect 547 633 560 635
rect 515 627 516 629
rect 518 627 519 629
rect 515 625 519 627
rect 575 629 579 658
rect 663 657 675 660
rect 647 654 659 655
rect 583 653 628 654
rect 583 651 584 653
rect 586 651 628 653
rect 583 650 628 651
rect 583 637 587 650
rect 624 646 628 650
rect 647 652 653 654
rect 655 652 659 654
rect 647 649 659 652
rect 647 647 649 649
rect 583 635 584 637
rect 586 635 587 637
rect 583 633 587 635
rect 591 642 620 646
rect 624 645 631 646
rect 624 643 627 645
rect 629 643 631 645
rect 624 642 631 643
rect 591 637 597 642
rect 616 639 620 642
rect 647 641 651 647
rect 663 645 667 647
rect 663 643 664 645
rect 666 643 667 645
rect 663 639 667 643
rect 591 635 594 637
rect 596 635 597 637
rect 591 633 597 635
rect 604 637 612 638
rect 604 635 606 637
rect 608 635 612 637
rect 604 634 612 635
rect 616 637 617 639
rect 619 638 620 639
rect 655 638 667 639
rect 619 637 628 638
rect 616 635 625 637
rect 627 635 628 637
rect 616 634 628 635
rect 655 636 660 638
rect 662 636 667 638
rect 607 630 612 634
rect 655 633 667 636
rect 607 629 620 630
rect 575 628 603 629
rect 575 626 577 628
rect 579 626 599 628
rect 601 626 603 628
rect 575 625 603 626
rect 607 627 617 629
rect 619 627 620 629
rect 607 625 620 627
rect 671 629 675 657
rect 666 628 675 629
rect 666 626 668 628
rect 670 626 675 628
rect 683 662 699 663
rect 683 660 695 662
rect 697 660 699 662
rect 683 658 699 660
rect 683 638 687 658
rect 731 665 743 671
rect 738 662 743 665
rect 738 660 740 662
rect 742 660 743 662
rect 683 636 684 638
rect 686 636 687 638
rect 683 630 687 636
rect 722 640 727 647
rect 738 653 743 660
rect 738 651 739 653
rect 741 651 743 653
rect 738 649 743 651
rect 722 638 723 640
rect 725 639 727 640
rect 725 638 735 639
rect 722 637 735 638
rect 722 635 732 637
rect 734 635 735 637
rect 722 633 735 635
rect 683 629 707 630
rect 683 627 703 629
rect 705 627 707 629
rect 683 626 707 627
rect 666 625 675 626
rect 76 619 252 620
rect 76 617 119 619
rect 121 617 133 619
rect 135 617 145 619
rect 147 617 163 619
rect 165 617 173 619
rect 175 617 243 619
rect 245 617 252 619
rect 76 612 252 617
rect 515 619 747 620
rect 515 617 518 619
rect 520 617 528 619
rect 530 617 588 619
rect 590 617 610 619
rect 612 617 626 619
rect 628 617 685 619
rect 687 617 738 619
rect 740 617 747 619
rect 515 612 747 617
rect 76 607 260 612
rect 76 605 83 607
rect 85 605 136 607
rect 138 605 207 607
rect 209 605 217 607
rect 219 605 237 607
rect 239 605 249 607
rect 251 605 260 607
rect 76 604 260 605
rect 487 607 747 612
rect 487 605 498 607
rect 500 605 542 607
rect 544 605 620 607
rect 622 605 630 607
rect 632 605 664 607
rect 666 605 674 607
rect 676 605 690 607
rect 692 605 702 607
rect 704 605 747 607
rect 487 604 747 605
rect 148 598 157 599
rect 116 597 140 598
rect 116 595 118 597
rect 120 595 140 597
rect 116 594 140 595
rect 88 590 101 591
rect 88 588 89 590
rect 91 588 101 590
rect 88 586 101 588
rect 88 585 98 586
rect 96 584 98 585
rect 100 584 101 586
rect 80 573 85 575
rect 80 571 82 573
rect 84 571 85 573
rect 80 567 85 571
rect 96 577 101 584
rect 136 589 140 594
rect 136 587 137 589
rect 139 587 140 589
rect 80 565 81 567
rect 83 565 85 567
rect 80 559 85 565
rect 80 553 92 559
rect 136 566 140 587
rect 124 564 140 566
rect 124 562 126 564
rect 128 562 130 564
rect 132 562 140 564
rect 124 561 140 562
rect 148 596 149 598
rect 151 596 153 598
rect 155 596 157 598
rect 148 595 157 596
rect 148 567 152 595
rect 156 589 168 591
rect 156 587 157 589
rect 159 587 168 589
rect 156 585 168 587
rect 193 590 198 591
rect 193 588 194 590
rect 196 588 198 590
rect 156 581 160 585
rect 156 579 157 581
rect 159 579 160 581
rect 156 577 160 579
rect 172 577 176 583
rect 193 582 198 588
rect 210 595 222 599
rect 210 593 218 595
rect 220 593 222 595
rect 193 581 207 582
rect 193 579 201 581
rect 203 579 207 581
rect 193 578 207 579
rect 174 575 176 577
rect 164 572 176 575
rect 164 570 166 572
rect 168 570 176 572
rect 164 569 176 570
rect 186 573 199 574
rect 186 571 191 573
rect 193 571 199 573
rect 186 570 199 571
rect 148 561 160 567
rect 186 564 190 570
rect 218 575 222 593
rect 218 573 219 575
rect 221 573 222 575
rect 186 562 187 564
rect 189 562 190 564
rect 186 561 190 562
rect 217 571 222 573
rect 217 569 218 571
rect 220 569 222 571
rect 217 564 222 569
rect 217 562 218 564
rect 220 562 222 564
rect 217 560 222 562
rect 234 590 238 599
rect 234 588 236 590
rect 234 572 238 588
rect 242 583 246 591
rect 499 597 511 599
rect 499 595 508 597
rect 510 595 511 597
rect 499 593 511 595
rect 529 598 559 599
rect 529 596 531 598
rect 533 596 553 598
rect 555 596 559 598
rect 529 594 559 596
rect 499 588 503 593
rect 516 589 541 590
rect 499 586 500 588
rect 502 586 503 588
rect 499 585 503 586
rect 507 586 511 588
rect 516 587 518 589
rect 520 587 523 589
rect 525 587 537 589
rect 539 587 541 589
rect 516 586 541 587
rect 547 587 551 589
rect 507 584 508 586
rect 510 584 511 586
rect 242 582 254 583
rect 242 581 247 582
rect 242 579 243 581
rect 245 580 247 581
rect 249 580 254 582
rect 507 582 511 584
rect 245 579 254 580
rect 242 577 254 579
rect 496 580 502 581
rect 496 578 498 580
rect 500 578 502 580
rect 507 578 520 582
rect 530 578 536 586
rect 547 585 548 587
rect 550 585 551 587
rect 496 574 502 578
rect 516 574 520 578
rect 547 574 551 585
rect 234 570 236 572
rect 234 567 238 570
rect 496 570 511 574
rect 516 573 551 574
rect 516 571 548 573
rect 550 571 551 573
rect 516 570 551 571
rect 234 565 246 567
rect 234 563 236 565
rect 238 563 239 565
rect 241 563 246 565
rect 234 561 246 563
rect 507 558 511 570
rect 555 566 559 594
rect 590 590 603 591
rect 590 588 591 590
rect 593 588 603 590
rect 590 585 603 588
rect 607 590 611 591
rect 607 588 608 590
rect 610 588 611 590
rect 563 580 567 582
rect 565 578 567 580
rect 590 581 596 585
rect 590 579 592 581
rect 594 579 596 581
rect 590 578 596 579
rect 607 582 611 588
rect 631 591 635 599
rect 633 589 635 591
rect 607 581 620 582
rect 607 579 614 581
rect 616 579 620 581
rect 607 578 620 579
rect 526 565 559 566
rect 526 563 528 565
rect 530 563 556 565
rect 558 563 559 565
rect 526 562 559 563
rect 563 558 567 578
rect 590 573 604 574
rect 590 571 600 573
rect 602 572 604 573
rect 606 572 612 574
rect 602 571 612 572
rect 590 570 612 571
rect 507 557 567 558
rect 507 555 564 557
rect 566 555 567 557
rect 507 554 567 555
rect 598 562 604 570
rect 631 570 635 589
rect 650 587 655 591
rect 650 585 652 587
rect 654 585 655 587
rect 667 595 679 599
rect 667 593 675 595
rect 677 593 679 595
rect 650 582 655 585
rect 650 581 664 582
rect 650 579 658 581
rect 660 579 664 581
rect 650 578 664 579
rect 633 568 635 570
rect 631 566 635 568
rect 622 565 635 566
rect 622 563 623 565
rect 625 563 635 565
rect 622 562 631 563
rect 630 561 631 562
rect 633 561 635 563
rect 643 573 656 574
rect 643 571 648 573
rect 650 571 653 573
rect 655 571 656 573
rect 643 570 656 571
rect 643 561 647 570
rect 675 573 679 593
rect 703 598 707 599
rect 703 596 704 598
rect 706 596 707 598
rect 695 583 699 591
rect 703 590 707 596
rect 734 598 743 599
rect 734 596 736 598
rect 738 596 743 598
rect 734 595 743 596
rect 705 588 707 590
rect 687 581 699 583
rect 687 580 696 581
rect 687 578 688 580
rect 690 579 696 580
rect 698 579 699 581
rect 690 578 699 579
rect 687 577 699 578
rect 674 571 679 573
rect 674 569 675 571
rect 677 569 679 571
rect 674 567 679 569
rect 703 572 707 588
rect 723 590 735 591
rect 723 588 724 590
rect 726 588 735 590
rect 723 585 735 588
rect 705 570 707 572
rect 703 567 707 570
rect 715 577 719 583
rect 731 581 735 585
rect 731 579 732 581
rect 734 579 735 581
rect 715 575 717 577
rect 731 577 735 579
rect 739 588 743 595
rect 739 586 740 588
rect 742 586 743 588
rect 715 572 727 575
rect 715 570 716 572
rect 718 570 727 572
rect 715 569 727 570
rect 739 567 743 586
rect 674 565 676 567
rect 678 565 679 567
rect 674 564 679 565
rect 630 553 635 561
rect 674 562 675 564
rect 677 562 679 564
rect 674 560 679 562
rect 695 565 707 567
rect 695 563 703 565
rect 705 563 707 565
rect 695 561 707 563
rect 731 561 743 567
rect 76 547 260 548
rect 76 545 116 547
rect 118 545 217 547
rect 219 545 237 547
rect 239 545 249 547
rect 251 545 260 547
rect 76 535 260 545
rect 487 547 747 548
rect 487 545 498 547
rect 500 545 520 547
rect 522 545 560 547
rect 562 545 586 547
rect 588 545 600 547
rect 602 545 674 547
rect 676 545 690 547
rect 692 545 702 547
rect 704 545 747 547
rect 487 540 747 545
rect 76 533 131 535
rect 133 533 143 535
rect 145 533 181 535
rect 183 533 233 535
rect 235 533 260 535
rect 76 532 260 533
rect 438 535 747 540
rect 438 533 448 535
rect 450 533 460 535
rect 462 533 480 535
rect 482 533 557 535
rect 559 533 634 535
rect 636 533 705 535
rect 707 533 747 535
rect 438 532 747 533
rect 96 518 102 520
rect 96 516 99 518
rect 101 516 102 518
rect 96 511 102 516
rect 136 517 148 519
rect 136 516 144 517
rect 136 514 139 516
rect 141 515 144 516
rect 146 515 148 517
rect 141 514 148 515
rect 136 513 148 514
rect 96 510 99 511
rect 80 509 99 510
rect 101 509 102 511
rect 80 507 81 509
rect 83 507 102 509
rect 80 506 102 507
rect 112 510 117 511
rect 112 508 114 510
rect 116 508 117 510
rect 80 486 84 506
rect 112 502 117 508
rect 144 510 148 513
rect 146 508 148 510
rect 100 501 117 502
rect 100 499 102 501
rect 104 499 117 501
rect 100 498 117 499
rect 128 501 140 503
rect 128 499 137 501
rect 139 499 140 501
rect 90 496 94 498
rect 128 497 140 499
rect 90 494 91 496
rect 93 494 94 496
rect 90 493 117 494
rect 90 491 91 493
rect 93 491 113 493
rect 115 491 117 493
rect 136 492 140 497
rect 90 490 117 491
rect 80 485 98 486
rect 80 483 91 485
rect 93 483 94 485
rect 96 483 98 485
rect 80 482 98 483
rect 112 481 117 490
rect 136 490 137 492
rect 139 490 140 492
rect 136 489 140 490
rect 144 492 148 508
rect 146 490 148 492
rect 144 481 148 490
rect 159 518 175 519
rect 159 516 171 518
rect 173 516 175 518
rect 159 514 175 516
rect 159 497 163 514
rect 207 526 219 527
rect 207 524 216 526
rect 218 524 219 526
rect 207 521 219 524
rect 198 502 203 503
rect 198 500 200 502
rect 202 500 203 502
rect 159 495 160 497
rect 162 495 163 497
rect 159 486 163 495
rect 198 496 203 500
rect 214 509 219 521
rect 453 518 465 519
rect 240 517 257 518
rect 240 515 242 517
rect 244 515 247 517
rect 249 515 257 517
rect 240 514 257 515
rect 214 507 215 509
rect 217 507 219 509
rect 214 505 219 507
rect 229 509 242 510
rect 229 507 239 509
rect 241 507 242 509
rect 229 506 242 507
rect 229 502 233 506
rect 198 494 199 496
rect 201 495 203 496
rect 201 494 211 495
rect 198 489 211 494
rect 229 500 231 502
rect 229 497 233 500
rect 253 495 257 514
rect 453 516 454 518
rect 456 517 465 518
rect 456 516 461 517
rect 453 515 461 516
rect 463 515 465 517
rect 453 513 465 515
rect 461 510 465 513
rect 463 508 465 510
rect 445 501 457 503
rect 445 500 454 501
rect 445 498 447 500
rect 449 499 454 500
rect 456 499 457 501
rect 449 498 457 499
rect 445 497 457 498
rect 237 492 257 495
rect 237 490 242 492
rect 244 490 257 492
rect 237 489 257 490
rect 453 489 457 497
rect 159 485 183 486
rect 159 483 179 485
rect 181 483 183 485
rect 461 492 465 508
rect 481 511 485 527
rect 489 525 494 527
rect 489 523 491 525
rect 493 523 494 525
rect 489 519 494 523
rect 489 518 525 519
rect 489 516 491 518
rect 493 516 511 518
rect 513 516 525 518
rect 489 515 525 516
rect 513 513 525 515
rect 481 510 493 511
rect 481 508 482 510
rect 484 508 493 510
rect 481 507 493 508
rect 463 490 465 492
rect 159 482 183 483
rect 461 481 465 490
rect 481 501 485 503
rect 481 499 482 501
rect 484 499 485 501
rect 481 495 485 499
rect 489 497 493 507
rect 503 508 509 511
rect 503 506 504 508
rect 506 506 509 508
rect 503 501 509 506
rect 497 497 509 501
rect 513 501 517 503
rect 513 499 514 501
rect 516 499 517 501
rect 513 498 517 499
rect 481 493 482 495
rect 484 493 485 495
rect 481 487 485 493
rect 497 492 501 497
rect 513 496 514 498
rect 516 496 517 498
rect 513 493 517 496
rect 497 490 498 492
rect 500 490 501 492
rect 481 481 493 487
rect 497 481 501 490
rect 505 489 517 493
rect 505 481 509 489
rect 521 485 525 513
rect 513 484 525 485
rect 513 482 515 484
rect 517 482 522 484
rect 524 482 525 484
rect 535 518 551 519
rect 535 516 547 518
rect 549 516 551 518
rect 535 514 551 516
rect 535 495 539 514
rect 583 526 595 527
rect 583 524 586 526
rect 588 524 595 526
rect 583 521 595 524
rect 535 493 536 495
rect 538 493 539 495
rect 535 486 539 493
rect 574 496 579 503
rect 590 509 595 521
rect 590 507 591 509
rect 593 507 595 509
rect 590 505 595 507
rect 603 518 607 519
rect 603 516 604 518
rect 606 516 607 518
rect 603 510 607 516
rect 666 525 672 526
rect 666 523 668 525
rect 670 523 672 525
rect 666 522 672 523
rect 666 520 667 522
rect 669 520 672 522
rect 634 518 639 520
rect 603 509 616 510
rect 603 507 608 509
rect 610 507 616 509
rect 603 506 616 507
rect 574 494 575 496
rect 577 495 579 496
rect 577 494 587 495
rect 574 492 587 494
rect 574 490 584 492
rect 586 490 587 492
rect 574 489 587 490
rect 610 501 624 502
rect 610 499 618 501
rect 620 499 624 501
rect 610 498 624 499
rect 634 516 635 518
rect 637 516 639 518
rect 634 511 639 516
rect 666 519 672 520
rect 666 518 675 519
rect 666 516 668 518
rect 670 516 675 518
rect 666 515 675 516
rect 634 509 635 511
rect 637 509 639 511
rect 634 507 639 509
rect 610 495 615 498
rect 610 493 611 495
rect 613 493 615 495
rect 610 489 615 493
rect 535 485 559 486
rect 535 483 555 485
rect 557 483 559 485
rect 635 487 639 507
rect 655 509 659 511
rect 655 507 656 509
rect 658 507 659 509
rect 655 503 667 507
rect 647 499 651 503
rect 663 501 667 503
rect 663 499 664 501
rect 666 499 667 501
rect 647 498 659 499
rect 647 496 654 498
rect 656 496 659 498
rect 663 497 667 499
rect 647 495 659 496
rect 655 492 659 495
rect 655 490 656 492
rect 658 490 659 492
rect 655 489 659 490
rect 535 482 559 483
rect 627 486 635 487
rect 627 484 628 486
rect 630 485 635 486
rect 637 485 639 487
rect 630 484 639 485
rect 513 481 525 482
rect 627 481 639 484
rect 671 487 675 515
rect 663 485 675 487
rect 658 484 675 485
rect 658 482 660 484
rect 662 482 675 484
rect 683 518 699 519
rect 683 517 695 518
rect 683 515 688 517
rect 690 516 695 517
rect 697 516 699 518
rect 690 515 699 516
rect 683 514 699 515
rect 683 492 687 514
rect 731 521 743 527
rect 738 516 743 521
rect 738 514 740 516
rect 742 514 743 516
rect 683 490 684 492
rect 686 490 687 492
rect 722 496 727 503
rect 738 509 743 514
rect 738 507 739 509
rect 741 507 743 509
rect 738 505 743 507
rect 722 494 723 496
rect 725 495 727 496
rect 725 494 735 495
rect 683 486 687 490
rect 722 493 735 494
rect 722 491 732 493
rect 734 491 735 493
rect 722 489 735 491
rect 683 485 707 486
rect 683 483 703 485
rect 705 483 707 485
rect 683 482 707 483
rect 658 481 675 482
rect 76 475 260 476
rect 76 473 119 475
rect 121 473 131 475
rect 133 473 143 475
rect 145 473 161 475
rect 163 473 214 475
rect 216 473 232 475
rect 234 473 252 475
rect 254 473 260 475
rect 76 468 260 473
rect 438 475 747 476
rect 438 473 448 475
rect 450 473 460 475
rect 462 473 483 475
rect 485 473 537 475
rect 539 473 590 475
rect 592 473 624 475
rect 626 473 634 475
rect 636 473 650 475
rect 652 473 671 475
rect 673 473 685 475
rect 687 473 738 475
rect 740 473 747 475
rect 438 468 747 473
rect 1 360 801 365
rect 1 358 8 360
rect 10 358 15 360
rect 17 358 108 360
rect 110 358 115 360
rect 117 358 208 360
rect 210 358 215 360
rect 217 358 308 360
rect 310 358 315 360
rect 317 358 408 360
rect 410 358 415 360
rect 417 358 508 360
rect 510 358 515 360
rect 517 358 608 360
rect 610 358 615 360
rect 617 358 708 360
rect 710 358 715 360
rect 717 358 801 360
rect 1 357 801 358
rect 77 351 81 357
rect 37 349 44 350
rect 37 347 40 349
rect 42 347 44 349
rect 37 346 44 347
rect 5 335 17 336
rect 5 333 6 335
rect 8 334 17 335
rect 8 333 12 334
rect 5 332 12 333
rect 14 332 17 334
rect 5 330 17 332
rect 5 325 9 330
rect 5 323 6 325
rect 8 323 9 325
rect 5 322 9 323
rect 37 325 41 346
rect 37 323 38 325
rect 40 323 41 325
rect 37 318 41 323
rect 37 316 38 318
rect 40 316 41 318
rect 37 311 41 316
rect 77 342 81 347
rect 77 340 78 342
rect 80 340 81 342
rect 77 336 81 340
rect 74 335 81 336
rect 74 333 76 335
rect 78 333 81 335
rect 85 341 89 351
rect 137 349 144 350
rect 137 347 140 349
rect 142 347 144 349
rect 137 346 144 347
rect 177 350 181 351
rect 177 348 178 350
rect 180 348 181 350
rect 85 339 86 341
rect 88 339 89 341
rect 85 337 89 339
rect 85 335 86 337
rect 88 335 89 337
rect 85 333 89 335
rect 74 332 81 333
rect 77 328 81 332
rect 77 322 89 328
rect 105 334 117 336
rect 105 332 112 334
rect 114 332 117 334
rect 105 330 117 332
rect 105 326 109 330
rect 105 324 106 326
rect 108 324 109 326
rect 105 323 109 324
rect 105 318 109 319
rect 105 316 107 318
rect 105 315 109 316
rect 137 325 141 346
rect 137 323 138 325
rect 140 323 141 325
rect 137 322 141 323
rect 137 320 138 322
rect 140 320 141 322
rect 137 318 141 320
rect 137 316 138 318
rect 140 316 141 318
rect 137 311 141 316
rect 177 336 181 348
rect 174 335 181 336
rect 174 333 176 335
rect 178 333 181 335
rect 185 341 189 351
rect 201 349 205 350
rect 185 339 186 341
rect 188 339 189 341
rect 185 337 189 339
rect 185 335 186 337
rect 188 335 189 337
rect 185 333 189 335
rect 174 332 181 333
rect 177 328 181 332
rect 177 322 189 328
rect 201 347 202 349
rect 204 347 205 349
rect 201 336 205 347
rect 237 349 244 350
rect 237 347 240 349
rect 242 347 244 349
rect 237 346 244 347
rect 277 349 281 350
rect 201 334 217 336
rect 201 332 212 334
rect 214 332 217 334
rect 205 330 217 332
rect 205 325 209 330
rect 205 323 206 325
rect 208 323 209 325
rect 205 322 209 323
rect 237 329 241 346
rect 237 327 238 329
rect 240 327 241 329
rect 237 325 241 327
rect 237 323 238 325
rect 240 323 241 325
rect 237 318 241 323
rect 237 316 238 318
rect 240 316 241 318
rect 237 311 241 316
rect 277 347 278 349
rect 280 347 281 349
rect 277 336 281 347
rect 274 335 281 336
rect 274 333 276 335
rect 278 333 281 335
rect 285 341 289 351
rect 337 349 344 350
rect 337 347 340 349
rect 342 347 344 349
rect 337 346 344 347
rect 285 339 286 341
rect 288 339 289 341
rect 285 337 289 339
rect 285 335 286 337
rect 288 335 289 337
rect 285 333 289 335
rect 274 332 281 333
rect 277 328 281 332
rect 277 322 289 328
rect 305 334 317 336
rect 305 333 312 334
rect 305 331 306 333
rect 308 332 312 333
rect 314 332 317 334
rect 308 331 317 332
rect 305 330 317 331
rect 305 326 309 330
rect 305 325 310 326
rect 305 323 307 325
rect 309 323 310 325
rect 305 322 310 323
rect 337 325 341 346
rect 337 323 338 325
rect 340 323 341 325
rect 337 318 341 323
rect 337 316 338 318
rect 340 316 341 318
rect 337 311 341 316
rect 376 347 389 351
rect 385 341 389 347
rect 437 349 444 350
rect 437 347 440 349
rect 442 347 444 349
rect 437 346 444 347
rect 385 339 386 341
rect 388 339 389 341
rect 385 337 389 339
rect 374 335 381 336
rect 374 333 376 335
rect 378 333 381 335
rect 385 335 386 337
rect 388 335 389 337
rect 385 333 389 335
rect 374 332 381 333
rect 377 328 381 332
rect 377 325 389 328
rect 377 323 386 325
rect 388 323 389 325
rect 377 322 389 323
rect 405 334 417 336
rect 405 332 412 334
rect 414 332 417 334
rect 405 330 417 332
rect 405 325 409 330
rect 405 323 406 325
rect 408 323 409 325
rect 405 322 409 323
rect 437 325 441 346
rect 437 323 438 325
rect 440 323 441 325
rect 437 321 441 323
rect 437 319 438 321
rect 440 319 441 321
rect 437 318 441 319
rect 437 316 438 318
rect 440 316 441 318
rect 437 311 441 316
rect 476 347 489 351
rect 500 349 504 350
rect 485 341 489 347
rect 485 339 486 341
rect 488 339 489 341
rect 485 337 489 339
rect 474 335 481 336
rect 474 333 476 335
rect 478 333 481 335
rect 485 335 486 337
rect 488 335 489 337
rect 485 333 489 335
rect 474 332 481 333
rect 477 331 481 332
rect 477 329 478 331
rect 480 329 481 331
rect 477 328 481 329
rect 477 322 489 328
rect 500 347 501 349
rect 503 347 504 349
rect 500 336 504 347
rect 537 349 544 350
rect 537 347 540 349
rect 542 347 544 349
rect 537 346 544 347
rect 500 334 517 336
rect 500 332 512 334
rect 514 332 517 334
rect 505 330 517 332
rect 505 322 509 330
rect 537 333 541 346
rect 537 331 538 333
rect 540 331 541 333
rect 537 325 541 331
rect 537 323 538 325
rect 540 323 541 325
rect 537 318 541 323
rect 537 316 538 318
rect 540 316 541 318
rect 537 311 541 316
rect 576 347 589 351
rect 600 350 604 351
rect 600 348 601 350
rect 603 348 604 350
rect 585 341 589 347
rect 585 339 586 341
rect 588 339 589 341
rect 585 337 589 339
rect 574 335 581 336
rect 574 333 576 335
rect 578 333 581 335
rect 585 335 586 337
rect 588 335 589 337
rect 585 333 589 335
rect 574 332 581 333
rect 577 328 581 332
rect 577 325 589 328
rect 577 323 586 325
rect 588 323 589 325
rect 577 322 589 323
rect 600 336 604 348
rect 637 349 644 350
rect 637 347 640 349
rect 642 347 644 349
rect 637 346 644 347
rect 600 334 617 336
rect 600 332 612 334
rect 614 332 617 334
rect 605 330 617 332
rect 605 328 609 330
rect 605 326 606 328
rect 608 326 609 328
rect 605 322 609 326
rect 637 333 641 346
rect 637 331 638 333
rect 640 331 641 333
rect 637 325 641 331
rect 637 323 638 325
rect 640 323 641 325
rect 637 318 641 323
rect 637 316 638 318
rect 640 316 641 318
rect 637 311 641 316
rect 676 347 689 351
rect 700 349 705 350
rect 685 341 689 347
rect 685 339 686 341
rect 688 339 689 341
rect 685 337 689 339
rect 674 335 681 336
rect 674 333 676 335
rect 678 333 681 335
rect 685 335 686 337
rect 688 335 689 337
rect 685 333 689 335
rect 674 332 681 333
rect 677 328 681 332
rect 677 325 689 328
rect 677 323 686 325
rect 688 323 689 325
rect 677 322 689 323
rect 700 347 702 349
rect 704 347 705 349
rect 700 336 705 347
rect 737 349 744 350
rect 737 347 740 349
rect 742 347 744 349
rect 737 346 744 347
rect 700 334 717 336
rect 700 332 712 334
rect 714 332 717 334
rect 705 330 717 332
rect 705 325 709 330
rect 705 323 706 325
rect 708 323 709 325
rect 705 322 709 323
rect 737 325 741 346
rect 737 323 738 325
rect 740 323 741 325
rect 737 318 741 323
rect 737 316 738 318
rect 740 316 741 318
rect 737 311 741 316
rect 776 347 789 351
rect 785 341 789 347
rect 785 339 786 341
rect 788 339 789 341
rect 785 337 789 339
rect 774 335 781 336
rect 774 333 776 335
rect 778 333 781 335
rect 785 335 786 337
rect 788 335 789 337
rect 785 333 789 335
rect 774 332 781 333
rect 777 328 781 332
rect 777 325 789 328
rect 777 323 786 325
rect 788 323 789 325
rect 777 322 789 323
rect 28 310 38 311
rect 28 308 29 310
rect 31 309 38 310
rect 40 309 41 311
rect 31 308 41 309
rect 28 307 41 308
rect 128 309 138 311
rect 140 309 141 311
rect 128 307 141 309
rect 228 309 238 311
rect 240 309 241 311
rect 228 307 241 309
rect 328 309 338 311
rect 340 309 341 311
rect 328 307 341 309
rect 428 309 438 311
rect 440 309 441 311
rect 428 307 441 309
rect 528 309 538 311
rect 540 309 541 311
rect 528 307 541 309
rect 628 309 638 311
rect 640 309 641 311
rect 628 307 641 309
rect 728 310 738 311
rect 728 308 729 310
rect 731 309 738 310
rect 740 309 741 311
rect 731 308 741 309
rect 728 307 741 308
rect 1 300 801 301
rect 1 298 8 300
rect 10 298 108 300
rect 110 298 208 300
rect 210 298 308 300
rect 310 298 408 300
rect 410 298 508 300
rect 510 298 608 300
rect 610 298 708 300
rect 710 298 801 300
rect 1 293 801 298
rect 1 288 803 293
rect 1 286 92 288
rect 94 286 192 288
rect 194 286 292 288
rect 294 286 392 288
rect 394 286 494 288
rect 496 286 594 288
rect 596 286 694 288
rect 696 286 794 288
rect 796 286 803 288
rect 1 285 803 286
rect 61 277 74 279
rect 61 275 62 277
rect 64 275 74 277
rect 161 277 174 279
rect 161 275 162 277
rect 164 275 174 277
rect 261 277 274 279
rect 261 275 262 277
rect 264 275 274 277
rect 361 277 374 279
rect 361 275 362 277
rect 364 275 374 277
rect 463 277 476 279
rect 463 275 464 277
rect 466 275 476 277
rect 563 277 576 279
rect 563 275 564 277
rect 566 275 576 277
rect 663 277 676 279
rect 663 275 664 277
rect 666 275 676 277
rect 763 277 776 279
rect 763 275 764 277
rect 766 275 776 277
rect 13 258 25 264
rect 21 256 25 258
rect 21 254 22 256
rect 24 254 25 256
rect 21 253 28 254
rect 13 251 17 253
rect 13 249 14 251
rect 16 249 17 251
rect 21 251 24 253
rect 26 251 28 253
rect 21 250 28 251
rect 13 247 17 249
rect 13 245 14 247
rect 16 245 17 247
rect 13 239 17 245
rect 13 235 26 239
rect 61 270 65 275
rect 61 268 62 270
rect 64 268 65 270
rect 61 263 65 268
rect 61 261 62 263
rect 64 261 65 263
rect 61 240 65 261
rect 93 256 97 264
rect 85 254 97 256
rect 85 252 88 254
rect 90 252 102 254
rect 85 250 102 252
rect 58 239 66 240
rect 58 237 60 239
rect 62 237 63 239
rect 65 237 66 239
rect 58 236 66 237
rect 98 239 102 250
rect 98 237 99 239
rect 101 237 102 239
rect 113 264 117 265
rect 113 262 114 264
rect 116 262 125 264
rect 113 258 125 262
rect 121 254 125 258
rect 121 253 128 254
rect 113 251 117 253
rect 113 249 114 251
rect 116 249 117 251
rect 121 251 124 253
rect 126 251 128 253
rect 121 250 128 251
rect 113 247 117 249
rect 113 245 114 247
rect 116 245 117 247
rect 113 239 117 245
rect 98 236 102 237
rect 113 235 126 239
rect 161 270 165 275
rect 161 268 162 270
rect 164 268 165 270
rect 161 263 165 268
rect 161 261 162 263
rect 164 261 165 263
rect 161 240 165 261
rect 193 263 202 264
rect 193 261 199 263
rect 201 261 202 263
rect 193 260 202 261
rect 193 257 197 260
rect 190 256 197 257
rect 185 254 191 256
rect 193 254 197 256
rect 185 252 188 254
rect 190 252 197 254
rect 185 250 197 252
rect 213 258 225 264
rect 221 256 225 258
rect 221 254 222 256
rect 224 254 225 256
rect 221 253 228 254
rect 213 251 217 253
rect 213 249 214 251
rect 216 249 217 251
rect 221 251 224 253
rect 226 251 228 253
rect 221 250 228 251
rect 213 247 217 249
rect 213 245 214 247
rect 216 245 217 247
rect 158 239 166 240
rect 158 237 160 239
rect 162 237 163 239
rect 165 237 166 239
rect 158 236 166 237
rect 213 239 217 245
rect 213 235 226 239
rect 261 270 265 275
rect 261 268 262 270
rect 264 268 265 270
rect 261 263 265 268
rect 261 261 262 263
rect 264 261 265 263
rect 261 240 265 261
rect 293 264 302 265
rect 293 262 299 264
rect 301 262 302 264
rect 293 261 302 262
rect 293 256 297 261
rect 285 254 297 256
rect 285 252 288 254
rect 290 252 297 254
rect 285 250 297 252
rect 313 264 317 265
rect 313 262 314 264
rect 316 262 325 264
rect 313 258 325 262
rect 321 254 325 258
rect 321 253 328 254
rect 313 251 317 253
rect 313 249 314 251
rect 316 249 317 251
rect 321 251 324 253
rect 326 251 328 253
rect 321 250 328 251
rect 313 247 317 249
rect 313 245 314 247
rect 316 245 317 247
rect 258 239 266 240
rect 258 237 260 239
rect 262 237 263 239
rect 265 237 266 239
rect 258 236 266 237
rect 313 239 317 245
rect 313 235 326 239
rect 361 270 365 275
rect 361 268 362 270
rect 364 268 365 270
rect 361 263 365 268
rect 361 261 362 263
rect 364 261 365 263
rect 361 240 365 261
rect 393 257 397 264
rect 390 256 397 257
rect 385 254 391 256
rect 393 254 397 256
rect 385 252 388 254
rect 390 252 404 254
rect 385 250 404 252
rect 358 239 366 240
rect 358 237 360 239
rect 362 237 363 239
rect 365 237 366 239
rect 358 236 366 237
rect 400 239 404 250
rect 400 237 401 239
rect 403 237 404 239
rect 415 258 427 264
rect 423 256 427 258
rect 423 254 424 256
rect 426 254 427 256
rect 423 253 430 254
rect 415 251 419 253
rect 415 249 416 251
rect 418 249 419 251
rect 423 251 426 253
rect 428 251 430 253
rect 423 250 430 251
rect 415 247 419 249
rect 415 245 416 247
rect 418 245 419 247
rect 415 239 419 245
rect 400 235 404 237
rect 415 235 428 239
rect 463 270 467 275
rect 463 268 464 270
rect 466 268 467 270
rect 463 263 467 268
rect 463 261 464 263
rect 466 261 467 263
rect 463 240 467 261
rect 495 264 504 265
rect 495 262 501 264
rect 503 262 504 264
rect 495 261 504 262
rect 495 256 499 261
rect 487 254 499 256
rect 487 252 490 254
rect 492 252 499 254
rect 487 250 499 252
rect 515 264 519 265
rect 515 262 516 264
rect 518 262 527 264
rect 515 258 527 262
rect 523 254 527 258
rect 523 253 530 254
rect 515 251 519 253
rect 515 249 516 251
rect 518 249 519 251
rect 523 251 526 253
rect 528 251 530 253
rect 523 250 530 251
rect 515 247 519 249
rect 515 245 516 247
rect 518 245 519 247
rect 460 239 468 240
rect 460 237 462 239
rect 464 237 465 239
rect 467 237 468 239
rect 460 236 468 237
rect 515 239 519 245
rect 515 235 528 239
rect 563 270 567 275
rect 563 268 564 270
rect 566 268 567 270
rect 563 263 567 268
rect 563 261 564 263
rect 566 261 567 263
rect 563 240 567 261
rect 595 257 599 264
rect 592 256 599 257
rect 587 254 593 256
rect 595 254 599 256
rect 587 252 590 254
rect 592 252 599 254
rect 587 250 599 252
rect 615 258 627 264
rect 623 256 627 258
rect 623 254 624 256
rect 626 254 627 256
rect 623 253 630 254
rect 615 251 619 253
rect 615 249 616 251
rect 618 249 619 251
rect 623 251 626 253
rect 628 251 630 253
rect 623 250 630 251
rect 615 247 619 249
rect 615 245 616 247
rect 618 245 619 247
rect 560 239 568 240
rect 560 237 562 239
rect 564 237 565 239
rect 567 237 568 239
rect 560 236 568 237
rect 615 239 619 245
rect 615 235 628 239
rect 663 270 667 275
rect 663 268 664 270
rect 666 268 667 270
rect 663 263 667 268
rect 663 261 664 263
rect 666 261 667 263
rect 663 240 667 261
rect 695 264 704 265
rect 695 262 701 264
rect 703 262 704 264
rect 695 261 704 262
rect 695 256 699 261
rect 687 254 699 256
rect 687 252 690 254
rect 692 252 699 254
rect 687 250 699 252
rect 715 264 719 265
rect 715 262 716 264
rect 718 262 727 264
rect 715 258 727 262
rect 723 254 727 258
rect 723 253 730 254
rect 715 251 719 253
rect 715 249 716 251
rect 718 249 719 251
rect 723 251 726 253
rect 728 251 730 253
rect 723 250 730 251
rect 715 247 719 249
rect 715 245 716 247
rect 718 245 719 247
rect 660 239 668 240
rect 660 237 662 239
rect 664 237 665 239
rect 667 237 668 239
rect 660 236 668 237
rect 715 239 719 245
rect 715 235 728 239
rect 763 270 767 275
rect 763 268 764 270
rect 766 268 767 270
rect 763 263 767 268
rect 763 261 764 263
rect 766 261 767 263
rect 763 240 767 261
rect 795 257 799 264
rect 792 256 799 257
rect 787 254 793 256
rect 795 254 799 256
rect 787 252 790 254
rect 792 252 799 254
rect 787 250 799 252
rect 760 239 768 240
rect 760 237 762 239
rect 764 237 765 239
rect 767 237 768 239
rect 760 236 768 237
rect 1 228 803 229
rect 1 226 85 228
rect 87 226 92 228
rect 94 226 185 228
rect 187 226 192 228
rect 194 226 285 228
rect 287 226 292 228
rect 294 226 385 228
rect 387 226 392 228
rect 394 226 487 228
rect 489 226 494 228
rect 496 226 587 228
rect 589 226 594 228
rect 596 226 687 228
rect 689 226 694 228
rect 696 226 787 228
rect 789 226 794 228
rect 796 226 803 228
rect 1 216 803 226
rect 1 214 85 216
rect 87 214 92 216
rect 94 214 185 216
rect 187 214 192 216
rect 194 214 285 216
rect 287 214 292 216
rect 294 214 385 216
rect 387 214 392 216
rect 394 214 487 216
rect 489 214 494 216
rect 496 214 587 216
rect 589 214 594 216
rect 596 214 687 216
rect 689 214 694 216
rect 696 214 787 216
rect 789 214 794 216
rect 796 214 803 216
rect 1 213 803 214
rect 13 203 26 207
rect 13 197 17 203
rect 13 195 14 197
rect 16 195 17 197
rect 13 193 17 195
rect 13 191 14 193
rect 16 191 17 193
rect 13 189 17 191
rect 21 191 28 192
rect 21 189 24 191
rect 26 189 28 191
rect 21 188 28 189
rect 58 205 65 206
rect 58 203 60 205
rect 62 203 65 205
rect 58 202 65 203
rect 98 205 102 206
rect 98 203 99 205
rect 101 203 102 205
rect 21 184 25 188
rect 13 181 25 184
rect 13 179 14 181
rect 16 179 25 181
rect 13 178 25 179
rect 61 181 65 202
rect 61 179 62 181
rect 64 179 65 181
rect 61 174 65 179
rect 61 172 62 174
rect 64 172 65 174
rect 61 171 65 172
rect 98 192 102 203
rect 85 190 102 192
rect 85 188 88 190
rect 90 188 102 190
rect 113 203 126 207
rect 85 186 97 188
rect 93 178 97 186
rect 113 197 117 203
rect 113 195 114 197
rect 116 195 117 197
rect 113 193 117 195
rect 113 191 114 193
rect 116 191 117 193
rect 113 189 117 191
rect 121 192 128 193
rect 121 190 124 192
rect 126 190 128 192
rect 121 189 128 190
rect 121 187 122 189
rect 124 188 128 189
rect 158 205 165 206
rect 158 203 160 205
rect 162 203 165 205
rect 158 202 165 203
rect 124 187 125 188
rect 121 184 125 187
rect 113 178 125 184
rect 61 169 62 171
rect 64 169 65 171
rect 161 181 165 202
rect 161 179 162 181
rect 164 179 165 181
rect 161 174 165 179
rect 161 172 162 174
rect 164 172 165 174
rect 61 167 65 169
rect 161 167 165 172
rect 213 203 226 207
rect 185 190 197 192
rect 185 188 188 190
rect 190 188 197 190
rect 185 186 197 188
rect 193 181 197 186
rect 193 179 194 181
rect 196 179 197 181
rect 193 178 197 179
rect 213 197 217 203
rect 213 195 214 197
rect 216 195 217 197
rect 213 193 217 195
rect 213 191 214 193
rect 216 191 217 193
rect 213 189 217 191
rect 221 191 228 192
rect 221 189 224 191
rect 226 189 228 191
rect 221 188 228 189
rect 258 205 265 206
rect 258 203 260 205
rect 262 203 265 205
rect 258 202 265 203
rect 297 206 301 207
rect 297 204 298 206
rect 300 204 301 206
rect 221 184 225 188
rect 213 181 225 184
rect 213 179 214 181
rect 216 179 225 181
rect 213 178 225 179
rect 261 181 265 202
rect 261 179 262 181
rect 264 179 265 181
rect 261 174 265 179
rect 261 172 262 174
rect 264 172 265 174
rect 261 167 265 172
rect 297 192 301 204
rect 285 190 301 192
rect 285 188 288 190
rect 290 189 301 190
rect 290 188 294 189
rect 285 187 294 188
rect 296 187 301 189
rect 285 186 301 187
rect 313 203 326 207
rect 293 178 297 186
rect 313 197 317 203
rect 313 195 314 197
rect 316 195 317 197
rect 313 193 317 195
rect 313 191 314 193
rect 316 191 317 193
rect 313 189 317 191
rect 321 192 328 194
rect 321 190 324 192
rect 326 190 328 192
rect 321 189 328 190
rect 321 187 322 189
rect 324 188 328 189
rect 358 205 365 206
rect 358 203 360 205
rect 362 203 365 205
rect 358 202 365 203
rect 392 208 402 209
rect 392 206 393 208
rect 395 206 402 208
rect 392 205 402 206
rect 324 187 325 188
rect 321 184 325 187
rect 313 178 325 184
rect 361 181 365 202
rect 361 179 362 181
rect 364 179 365 181
rect 361 174 365 179
rect 361 172 362 174
rect 364 172 365 174
rect 361 167 365 172
rect 398 192 402 205
rect 385 190 402 192
rect 385 188 387 190
rect 389 188 402 190
rect 385 187 402 188
rect 415 203 428 207
rect 385 186 396 187
rect 392 181 396 186
rect 392 179 393 181
rect 395 179 396 181
rect 392 178 396 179
rect 415 197 419 203
rect 415 195 416 197
rect 418 195 419 197
rect 415 193 419 195
rect 415 191 416 193
rect 418 191 419 193
rect 415 189 419 191
rect 423 191 430 192
rect 423 189 426 191
rect 428 189 430 191
rect 423 188 430 189
rect 460 205 467 206
rect 460 203 462 205
rect 464 203 467 205
rect 460 202 467 203
rect 423 184 427 188
rect 415 181 427 184
rect 415 179 416 181
rect 418 179 427 181
rect 415 178 427 179
rect 463 181 467 202
rect 463 179 464 181
rect 466 179 467 181
rect 463 174 467 179
rect 463 172 464 174
rect 466 172 467 174
rect 463 167 467 172
rect 515 203 528 207
rect 487 190 499 192
rect 487 188 490 190
rect 492 189 499 190
rect 492 188 496 189
rect 487 187 496 188
rect 498 187 499 189
rect 487 186 499 187
rect 495 178 499 186
rect 515 197 519 203
rect 515 195 516 197
rect 518 195 519 197
rect 515 193 519 195
rect 515 191 516 193
rect 518 191 519 193
rect 515 189 519 191
rect 523 192 530 193
rect 523 190 526 192
rect 528 190 530 192
rect 523 189 530 190
rect 523 187 524 189
rect 526 188 530 189
rect 560 205 567 206
rect 560 203 562 205
rect 564 203 567 205
rect 560 202 567 203
rect 526 187 527 188
rect 523 184 527 187
rect 515 178 527 184
rect 563 181 567 202
rect 563 179 564 181
rect 566 179 567 181
rect 563 174 567 179
rect 563 172 564 174
rect 566 172 567 174
rect 563 167 567 172
rect 615 203 628 207
rect 587 190 599 192
rect 587 188 590 190
rect 592 188 599 190
rect 587 186 599 188
rect 595 181 599 186
rect 595 179 596 181
rect 598 179 599 181
rect 595 178 599 179
rect 615 197 619 203
rect 615 195 616 197
rect 618 195 619 197
rect 615 193 619 195
rect 615 191 616 193
rect 618 191 619 193
rect 615 189 619 191
rect 623 191 630 192
rect 623 189 626 191
rect 628 189 630 191
rect 623 188 630 189
rect 660 205 667 206
rect 660 203 662 205
rect 664 203 667 205
rect 660 202 667 203
rect 623 184 627 188
rect 615 181 627 184
rect 615 179 616 181
rect 618 179 627 181
rect 615 178 627 179
rect 663 181 667 202
rect 663 179 664 181
rect 666 179 667 181
rect 663 174 667 179
rect 663 172 664 174
rect 666 172 667 174
rect 663 167 667 172
rect 715 203 728 207
rect 687 190 699 192
rect 687 188 690 190
rect 692 189 699 190
rect 692 188 696 189
rect 687 187 696 188
rect 698 187 699 189
rect 687 186 699 187
rect 695 178 699 186
rect 715 197 719 203
rect 715 195 716 197
rect 718 195 719 197
rect 715 193 719 195
rect 715 191 716 193
rect 718 191 719 193
rect 715 189 719 191
rect 723 192 730 193
rect 723 190 726 192
rect 728 190 730 192
rect 723 189 730 190
rect 723 187 724 189
rect 726 188 730 189
rect 760 205 767 206
rect 760 203 762 205
rect 764 203 767 205
rect 760 202 767 203
rect 726 187 727 188
rect 723 184 727 187
rect 715 178 727 184
rect 763 181 767 202
rect 763 179 764 181
rect 766 179 767 181
rect 763 174 767 179
rect 763 172 764 174
rect 766 172 767 174
rect 763 167 767 172
rect 787 191 814 192
rect 787 190 811 191
rect 787 188 790 190
rect 792 189 811 190
rect 813 189 814 191
rect 792 188 814 189
rect 787 186 799 188
rect 795 182 799 186
rect 794 181 799 182
rect 794 179 795 181
rect 797 179 799 181
rect 794 178 799 179
rect 61 165 62 167
rect 64 165 74 167
rect 61 163 74 165
rect 161 165 162 167
rect 164 166 174 167
rect 164 165 171 166
rect 161 164 171 165
rect 173 164 174 166
rect 161 163 174 164
rect 261 165 262 167
rect 264 166 274 167
rect 264 165 271 166
rect 261 164 271 165
rect 273 164 274 166
rect 261 163 274 164
rect 361 165 362 167
rect 364 166 374 167
rect 364 165 371 166
rect 361 164 371 165
rect 373 164 374 166
rect 361 163 374 164
rect 463 165 464 167
rect 466 166 476 167
rect 466 165 473 166
rect 463 164 473 165
rect 475 164 476 166
rect 463 163 476 164
rect 563 165 564 167
rect 566 166 576 167
rect 566 165 573 166
rect 563 164 573 165
rect 575 164 576 166
rect 563 163 576 164
rect 663 165 664 167
rect 666 166 676 167
rect 666 165 673 166
rect 663 164 673 165
rect 675 164 676 166
rect 663 163 676 164
rect 763 165 764 167
rect 766 166 776 167
rect 766 165 773 166
rect 763 164 773 165
rect 775 164 776 166
rect 763 163 776 164
rect 1 156 803 157
rect 1 154 92 156
rect 94 154 192 156
rect 194 154 292 156
rect 294 154 392 156
rect 394 154 494 156
rect 496 154 594 156
rect 596 154 694 156
rect 696 154 794 156
rect 796 154 803 156
rect 1 144 803 154
rect 1 142 92 144
rect 94 142 192 144
rect 194 142 292 144
rect 294 142 392 144
rect 394 142 494 144
rect 496 142 594 144
rect 596 142 694 144
rect 696 142 794 144
rect 796 142 803 144
rect 1 141 803 142
rect 61 133 74 135
rect 61 131 62 133
rect 64 131 74 133
rect 161 133 174 135
rect 161 131 162 133
rect 164 131 174 133
rect 261 133 274 135
rect 261 131 262 133
rect 264 131 274 133
rect 361 133 374 135
rect 361 131 362 133
rect 364 131 374 133
rect 463 133 476 135
rect 463 131 464 133
rect 466 131 476 133
rect 563 133 576 135
rect 563 131 564 133
rect 566 131 576 133
rect 663 133 676 135
rect 663 131 664 133
rect 666 131 676 133
rect 763 133 776 135
rect 763 131 764 133
rect 766 131 776 133
rect 13 119 25 120
rect 13 117 14 119
rect 16 117 25 119
rect 13 114 25 117
rect 21 110 25 114
rect 21 109 28 110
rect 13 107 17 109
rect 13 105 14 107
rect 16 105 17 107
rect 21 107 24 109
rect 26 107 28 109
rect 21 106 28 107
rect 13 95 17 105
rect 13 94 26 95
rect 61 126 65 131
rect 61 124 62 126
rect 64 124 65 126
rect 61 119 65 124
rect 61 117 62 119
rect 64 117 65 119
rect 61 115 65 117
rect 61 113 62 115
rect 64 113 65 115
rect 61 96 65 113
rect 93 119 97 120
rect 93 117 94 119
rect 96 117 97 119
rect 93 112 97 117
rect 85 110 97 112
rect 85 108 88 110
rect 90 108 97 110
rect 85 106 97 108
rect 113 117 125 121
rect 121 112 125 117
rect 121 111 128 112
rect 121 109 122 111
rect 124 109 128 111
rect 113 107 117 109
rect 113 105 114 107
rect 116 105 117 107
rect 121 107 125 109
rect 127 107 128 109
rect 121 106 128 107
rect 13 92 23 94
rect 25 92 26 94
rect 13 91 26 92
rect 58 95 65 96
rect 58 93 60 95
rect 62 93 65 95
rect 58 92 65 93
rect 113 95 117 105
rect 113 94 126 95
rect 161 126 165 131
rect 261 130 265 131
rect 261 128 262 130
rect 264 128 265 130
rect 161 124 162 126
rect 164 124 165 126
rect 161 119 165 124
rect 161 117 162 119
rect 164 117 165 119
rect 161 103 165 117
rect 161 101 162 103
rect 164 101 165 103
rect 161 96 165 101
rect 193 119 201 120
rect 193 117 198 119
rect 200 117 201 119
rect 193 116 201 117
rect 193 112 197 116
rect 185 110 197 112
rect 185 108 188 110
rect 190 108 197 110
rect 185 106 197 108
rect 213 114 225 120
rect 221 110 225 114
rect 221 109 228 110
rect 213 107 217 109
rect 213 105 214 107
rect 216 105 217 107
rect 113 92 122 94
rect 124 92 126 94
rect 113 91 126 92
rect 158 95 165 96
rect 158 93 160 95
rect 162 93 165 95
rect 158 92 165 93
rect 213 95 217 105
rect 221 107 224 109
rect 226 107 228 109
rect 221 103 228 107
rect 221 101 222 103
rect 224 101 225 103
rect 221 100 225 101
rect 213 94 226 95
rect 261 126 265 128
rect 261 124 262 126
rect 264 124 265 126
rect 261 119 265 124
rect 261 117 262 119
rect 264 117 265 119
rect 261 96 265 117
rect 293 119 297 120
rect 293 117 294 119
rect 296 117 297 119
rect 293 112 297 117
rect 285 111 297 112
rect 285 110 294 111
rect 285 108 288 110
rect 290 109 294 110
rect 296 109 297 111
rect 290 108 297 109
rect 285 106 297 108
rect 313 119 325 120
rect 313 117 314 119
rect 316 117 325 119
rect 313 114 325 117
rect 321 110 325 114
rect 321 109 328 110
rect 313 107 317 109
rect 313 105 314 107
rect 316 105 317 107
rect 321 107 324 109
rect 326 107 328 109
rect 321 106 328 107
rect 213 92 222 94
rect 224 92 226 94
rect 213 91 226 92
rect 258 95 265 96
rect 258 93 260 95
rect 262 93 265 95
rect 258 92 265 93
rect 313 95 317 105
rect 313 94 326 95
rect 361 126 365 131
rect 361 124 362 126
rect 364 124 365 126
rect 361 119 365 124
rect 361 117 362 119
rect 364 117 365 119
rect 361 111 365 117
rect 361 109 362 111
rect 364 109 365 111
rect 361 96 365 109
rect 393 119 397 120
rect 393 117 394 119
rect 396 117 397 119
rect 393 112 397 117
rect 385 110 397 112
rect 385 108 388 110
rect 390 108 397 110
rect 385 106 397 108
rect 415 119 427 120
rect 415 117 416 119
rect 418 117 427 119
rect 415 114 427 117
rect 423 110 427 114
rect 423 109 430 110
rect 415 107 419 109
rect 415 105 416 107
rect 418 105 419 107
rect 423 107 426 109
rect 428 107 430 109
rect 423 106 430 107
rect 313 92 322 94
rect 324 92 326 94
rect 313 91 326 92
rect 358 95 365 96
rect 358 93 360 95
rect 362 93 365 95
rect 358 92 365 93
rect 415 95 419 105
rect 415 94 428 95
rect 463 126 467 131
rect 563 130 567 131
rect 563 128 564 130
rect 566 128 567 130
rect 663 130 667 131
rect 663 128 664 130
rect 666 128 667 130
rect 463 124 464 126
rect 466 124 467 126
rect 463 123 467 124
rect 463 121 464 123
rect 466 121 467 123
rect 463 119 467 121
rect 463 117 464 119
rect 466 117 467 119
rect 463 96 467 117
rect 495 119 499 120
rect 495 117 496 119
rect 498 117 499 119
rect 495 112 499 117
rect 487 110 499 112
rect 487 108 490 110
rect 492 108 499 110
rect 487 106 499 108
rect 515 114 527 120
rect 523 112 527 114
rect 523 110 524 112
rect 526 110 527 112
rect 523 109 530 110
rect 515 107 519 109
rect 515 105 516 107
rect 518 105 519 107
rect 523 107 526 109
rect 528 107 530 109
rect 523 106 530 107
rect 415 92 424 94
rect 426 92 428 94
rect 415 91 428 92
rect 460 95 467 96
rect 460 93 462 95
rect 464 93 467 95
rect 460 92 467 93
rect 515 95 519 105
rect 515 94 528 95
rect 563 126 567 128
rect 563 124 564 126
rect 566 124 567 126
rect 563 119 567 124
rect 563 117 564 119
rect 566 117 567 119
rect 563 96 567 117
rect 595 112 599 120
rect 587 110 599 112
rect 587 108 590 110
rect 592 108 603 110
rect 587 106 603 108
rect 599 103 603 106
rect 599 101 600 103
rect 602 101 603 103
rect 599 100 603 101
rect 615 120 619 121
rect 615 118 616 120
rect 618 118 627 120
rect 615 114 627 118
rect 623 110 627 114
rect 623 109 630 110
rect 615 107 619 109
rect 615 105 616 107
rect 618 105 619 107
rect 623 107 626 109
rect 628 107 630 109
rect 623 106 630 107
rect 515 92 525 94
rect 527 92 528 94
rect 515 91 528 92
rect 560 95 567 96
rect 560 93 562 95
rect 564 93 567 95
rect 560 92 567 93
rect 615 95 619 105
rect 615 94 628 95
rect 663 126 667 128
rect 663 124 664 126
rect 666 124 667 126
rect 663 119 667 124
rect 663 117 664 119
rect 666 117 667 119
rect 663 96 667 117
rect 695 119 704 120
rect 695 117 701 119
rect 703 117 704 119
rect 695 115 704 117
rect 695 113 699 115
rect 692 112 699 113
rect 687 110 693 112
rect 695 110 699 112
rect 687 108 690 110
rect 692 108 699 110
rect 687 106 699 108
rect 715 114 727 120
rect 723 110 727 114
rect 723 109 730 110
rect 715 107 719 109
rect 715 105 716 107
rect 718 105 719 107
rect 615 92 625 94
rect 627 92 628 94
rect 615 91 628 92
rect 660 95 667 96
rect 660 93 662 95
rect 664 93 667 95
rect 660 92 667 93
rect 715 95 719 105
rect 723 107 726 109
rect 728 107 730 109
rect 723 106 730 107
rect 723 104 724 106
rect 726 104 730 106
rect 723 103 730 104
rect 715 94 728 95
rect 763 126 767 131
rect 763 124 764 126
rect 766 124 767 126
rect 763 119 767 124
rect 763 117 764 119
rect 766 117 767 119
rect 763 98 767 117
rect 763 96 764 98
rect 766 96 767 98
rect 794 119 814 120
rect 794 117 795 119
rect 797 117 811 119
rect 813 117 814 119
rect 794 116 814 117
rect 795 112 799 116
rect 787 110 799 112
rect 787 108 790 110
rect 792 108 799 110
rect 787 106 799 108
rect 715 92 725 94
rect 727 92 728 94
rect 715 91 728 92
rect 760 95 767 96
rect 760 93 762 95
rect 764 93 767 95
rect 760 92 767 93
rect 1 84 803 85
rect 1 82 85 84
rect 87 82 92 84
rect 94 82 185 84
rect 187 82 192 84
rect 194 82 285 84
rect 287 82 292 84
rect 294 82 385 84
rect 387 82 392 84
rect 394 82 487 84
rect 489 82 494 84
rect 496 82 587 84
rect 589 82 594 84
rect 596 82 687 84
rect 689 82 694 84
rect 696 82 787 84
rect 789 82 794 84
rect 796 82 803 84
rect 1 77 803 82
rect 1 72 801 77
rect 1 70 8 72
rect 10 70 15 72
rect 17 70 108 72
rect 110 70 115 72
rect 117 70 208 72
rect 210 70 215 72
rect 217 70 308 72
rect 310 70 315 72
rect 317 70 408 72
rect 410 70 415 72
rect 417 70 508 72
rect 510 70 515 72
rect 517 70 608 72
rect 610 70 615 72
rect 617 70 708 72
rect 710 70 715 72
rect 717 70 801 72
rect 1 69 801 70
rect 77 63 81 69
rect 37 61 44 62
rect 37 59 40 61
rect 42 59 44 61
rect 37 58 44 59
rect 5 46 17 48
rect 5 44 12 46
rect 14 44 17 46
rect 5 42 17 44
rect 5 37 9 42
rect 5 35 6 37
rect 8 35 9 37
rect 5 34 9 35
rect 37 37 41 58
rect 37 35 38 37
rect 40 35 41 37
rect 37 30 41 35
rect 37 28 38 30
rect 40 28 41 30
rect 37 23 41 28
rect 77 54 81 59
rect 77 52 78 54
rect 80 52 81 54
rect 77 48 81 52
rect 74 47 81 48
rect 74 45 76 47
rect 78 45 81 47
rect 85 53 89 63
rect 137 61 144 62
rect 137 59 140 61
rect 142 59 144 61
rect 137 58 144 59
rect 177 62 181 63
rect 177 60 178 62
rect 180 60 181 62
rect 85 51 86 53
rect 88 51 89 53
rect 85 49 89 51
rect 85 47 86 49
rect 88 47 89 49
rect 85 45 89 47
rect 74 44 81 45
rect 77 40 81 44
rect 77 34 89 40
rect 105 46 117 48
rect 105 44 112 46
rect 114 44 117 46
rect 105 42 117 44
rect 105 38 109 42
rect 105 36 106 38
rect 108 36 109 38
rect 105 35 109 36
rect 105 30 109 31
rect 105 28 107 30
rect 105 27 109 28
rect 137 44 141 58
rect 137 42 138 44
rect 140 42 141 44
rect 137 37 141 42
rect 137 35 138 37
rect 140 35 141 37
rect 137 30 141 35
rect 137 28 138 30
rect 140 28 141 30
rect 137 23 141 28
rect 177 48 181 60
rect 174 47 181 48
rect 174 45 176 47
rect 178 45 181 47
rect 185 53 189 63
rect 237 61 244 62
rect 237 59 240 61
rect 242 59 244 61
rect 237 58 244 59
rect 277 61 281 62
rect 185 51 186 53
rect 188 51 189 53
rect 185 49 189 51
rect 185 47 186 49
rect 188 47 189 49
rect 185 45 189 47
rect 174 44 181 45
rect 177 40 181 44
rect 177 34 189 40
rect 205 46 217 48
rect 205 44 212 46
rect 214 44 217 46
rect 205 42 217 44
rect 205 37 209 42
rect 205 35 206 37
rect 208 35 209 37
rect 205 34 209 35
rect 237 41 241 58
rect 237 39 238 41
rect 240 39 241 41
rect 237 37 241 39
rect 237 35 238 37
rect 240 35 241 37
rect 237 30 241 35
rect 237 28 238 30
rect 240 28 241 30
rect 237 23 241 28
rect 277 59 278 61
rect 280 59 281 61
rect 277 48 281 59
rect 274 47 281 48
rect 274 45 276 47
rect 278 45 281 47
rect 285 53 289 63
rect 337 61 344 62
rect 337 59 340 61
rect 342 59 344 61
rect 337 58 344 59
rect 285 51 286 53
rect 288 51 289 53
rect 285 49 289 51
rect 285 47 286 49
rect 288 47 289 49
rect 285 45 289 47
rect 274 44 281 45
rect 277 40 281 44
rect 277 34 289 40
rect 305 46 317 48
rect 305 45 312 46
rect 305 43 306 45
rect 308 44 312 45
rect 314 44 317 46
rect 308 43 317 44
rect 305 42 317 43
rect 305 34 309 42
rect 337 37 341 58
rect 337 35 338 37
rect 340 35 341 37
rect 337 34 341 35
rect 337 32 338 34
rect 340 32 341 34
rect 337 30 341 32
rect 337 28 338 30
rect 340 28 341 30
rect 337 23 341 28
rect 376 59 389 63
rect 385 53 389 59
rect 437 61 444 62
rect 437 59 440 61
rect 442 59 444 61
rect 437 58 444 59
rect 385 51 386 53
rect 388 51 389 53
rect 385 49 389 51
rect 374 47 381 48
rect 374 45 376 47
rect 378 45 381 47
rect 385 47 386 49
rect 388 47 389 49
rect 385 45 389 47
rect 374 44 381 45
rect 377 40 381 44
rect 377 37 389 40
rect 377 35 386 37
rect 388 35 389 37
rect 377 34 389 35
rect 405 46 417 48
rect 405 44 412 46
rect 414 44 417 46
rect 405 42 417 44
rect 405 37 409 42
rect 405 35 406 37
rect 408 35 409 37
rect 405 34 409 35
rect 437 37 441 58
rect 437 35 438 37
rect 440 35 441 37
rect 437 33 441 35
rect 437 31 438 33
rect 440 31 441 33
rect 437 30 441 31
rect 437 28 438 30
rect 440 28 441 30
rect 437 23 441 28
rect 476 59 489 63
rect 500 61 504 62
rect 485 53 489 59
rect 485 51 486 53
rect 488 51 489 53
rect 485 49 489 51
rect 474 47 481 48
rect 474 45 476 47
rect 478 45 481 47
rect 485 47 486 49
rect 488 47 489 49
rect 485 45 489 47
rect 474 44 481 45
rect 477 43 481 44
rect 477 41 478 43
rect 480 41 481 43
rect 477 40 481 41
rect 477 34 489 40
rect 500 59 501 61
rect 503 59 504 61
rect 500 48 504 59
rect 537 61 544 62
rect 537 59 540 61
rect 542 59 544 61
rect 537 58 544 59
rect 500 46 517 48
rect 500 45 512 46
rect 500 44 506 45
rect 505 43 506 44
rect 508 44 512 45
rect 514 44 517 46
rect 508 43 517 44
rect 505 42 517 43
rect 505 34 509 42
rect 537 37 541 58
rect 537 35 538 37
rect 540 35 541 37
rect 537 33 541 35
rect 537 31 538 33
rect 540 31 541 33
rect 537 30 541 31
rect 537 28 538 30
rect 540 28 541 30
rect 537 23 541 28
rect 576 59 589 63
rect 600 62 604 63
rect 600 60 601 62
rect 603 60 604 62
rect 585 53 589 59
rect 585 51 586 53
rect 588 51 589 53
rect 585 49 589 51
rect 574 47 581 48
rect 574 45 576 47
rect 578 45 581 47
rect 585 47 586 49
rect 588 47 589 49
rect 585 45 589 47
rect 574 44 581 45
rect 577 40 581 44
rect 577 37 589 40
rect 577 35 586 37
rect 588 35 589 37
rect 577 34 589 35
rect 600 48 604 60
rect 637 61 644 62
rect 637 59 640 61
rect 642 59 644 61
rect 637 58 644 59
rect 600 46 617 48
rect 600 44 612 46
rect 614 44 617 46
rect 605 42 617 44
rect 605 34 609 42
rect 637 37 641 58
rect 637 35 638 37
rect 640 35 641 37
rect 637 30 641 35
rect 637 28 638 30
rect 640 28 641 30
rect 637 27 641 28
rect 637 25 638 27
rect 640 25 641 27
rect 676 59 689 63
rect 700 61 705 62
rect 685 53 689 59
rect 685 51 686 53
rect 688 51 689 53
rect 685 49 689 51
rect 674 47 681 48
rect 674 45 676 47
rect 678 45 681 47
rect 685 47 686 49
rect 688 47 689 49
rect 685 45 689 47
rect 674 44 681 45
rect 677 40 681 44
rect 677 37 689 40
rect 677 35 686 37
rect 688 35 689 37
rect 677 34 689 35
rect 700 59 702 61
rect 704 59 705 61
rect 700 48 705 59
rect 737 61 744 62
rect 737 59 740 61
rect 742 59 744 61
rect 737 58 744 59
rect 700 46 717 48
rect 700 44 712 46
rect 714 44 717 46
rect 705 42 717 44
rect 705 34 709 42
rect 737 37 741 58
rect 737 35 738 37
rect 740 35 741 37
rect 737 33 741 35
rect 737 31 738 33
rect 740 31 741 33
rect 737 30 741 31
rect 737 28 738 30
rect 740 28 741 30
rect 637 23 641 25
rect 737 23 741 28
rect 776 59 789 63
rect 785 53 789 59
rect 785 51 786 53
rect 788 51 789 53
rect 785 49 789 51
rect 774 47 781 48
rect 774 45 776 47
rect 778 45 781 47
rect 785 47 786 49
rect 788 47 789 49
rect 785 45 789 47
rect 774 44 781 45
rect 777 40 781 44
rect 777 37 789 40
rect 777 35 786 37
rect 788 35 789 37
rect 777 34 789 35
rect 28 22 38 23
rect 28 20 29 22
rect 31 21 38 22
rect 40 21 41 23
rect 31 20 41 21
rect 28 19 41 20
rect 128 21 138 23
rect 140 21 141 23
rect 128 19 141 21
rect 228 21 238 23
rect 240 21 241 23
rect 228 19 241 21
rect 328 21 338 23
rect 340 21 341 23
rect 328 19 341 21
rect 428 21 438 23
rect 440 21 441 23
rect 428 19 441 21
rect 528 21 538 23
rect 540 21 541 23
rect 528 19 541 21
rect 628 21 638 23
rect 640 21 641 23
rect 628 19 641 21
rect 728 21 738 23
rect 740 21 741 23
rect 728 19 741 21
rect 1 12 801 13
rect 1 10 8 12
rect 10 10 108 12
rect 110 10 208 12
rect 210 10 308 12
rect 310 10 408 12
rect 410 10 508 12
rect 510 10 608 12
rect 610 10 708 12
rect 710 10 801 12
rect 1 5 801 10
rect -16 -28 932 -23
rect -16 -30 -9 -28
rect -7 -30 97 -28
rect 99 -30 203 -28
rect 205 -30 309 -28
rect 311 -30 415 -28
rect 417 -30 521 -28
rect 523 -30 627 -28
rect 629 -30 733 -28
rect 735 -30 839 -28
rect 841 -30 932 -28
rect -16 -31 932 -30
rect 11 -39 24 -37
rect 11 -41 21 -39
rect 23 -41 24 -39
rect 117 -39 130 -37
rect 117 -41 127 -39
rect 129 -41 130 -39
rect 223 -39 236 -37
rect 223 -41 233 -39
rect 235 -41 236 -39
rect 329 -39 342 -37
rect 329 -41 339 -39
rect 341 -41 342 -39
rect 435 -39 448 -37
rect 435 -41 445 -39
rect 447 -41 448 -39
rect 541 -39 554 -37
rect 541 -41 551 -39
rect 553 -41 554 -39
rect 647 -39 660 -37
rect 647 -41 657 -39
rect 659 -41 660 -39
rect 753 -39 766 -37
rect 753 -41 763 -39
rect 765 -41 766 -39
rect 859 -39 872 -37
rect 859 -41 869 -39
rect 871 -41 872 -39
rect -12 -60 -8 -52
rect -12 -62 0 -60
rect -12 -64 -11 -62
rect -9 -64 -5 -62
rect -3 -64 0 -62
rect -12 -66 0 -64
rect 20 -46 24 -41
rect 20 -48 21 -46
rect 23 -48 24 -46
rect 20 -53 24 -48
rect 20 -55 21 -53
rect 23 -55 24 -53
rect 20 -76 24 -55
rect 60 -54 72 -52
rect 60 -56 68 -54
rect 70 -56 72 -54
rect 60 -58 72 -56
rect 60 -62 64 -58
rect 20 -77 27 -76
rect 20 -79 23 -77
rect 25 -79 27 -77
rect 20 -80 27 -79
rect 57 -63 64 -62
rect 57 -65 59 -63
rect 61 -65 64 -63
rect 57 -66 64 -65
rect 68 -65 72 -63
rect 68 -67 69 -65
rect 71 -67 72 -65
rect 68 -77 72 -67
rect 94 -53 98 -52
rect 94 -55 95 -53
rect 97 -55 98 -53
rect 94 -60 98 -55
rect 94 -62 106 -60
rect 94 -64 101 -62
rect 103 -64 106 -62
rect 94 -66 106 -64
rect 59 -78 72 -77
rect 126 -46 130 -41
rect 126 -48 127 -46
rect 129 -48 130 -46
rect 126 -53 130 -48
rect 126 -55 127 -53
rect 129 -55 130 -53
rect 126 -76 130 -55
rect 166 -54 178 -52
rect 166 -56 174 -54
rect 176 -56 178 -54
rect 166 -58 178 -56
rect 166 -62 170 -58
rect 59 -80 61 -78
rect 63 -80 72 -78
rect 59 -81 72 -80
rect 126 -77 133 -76
rect 126 -79 129 -77
rect 131 -79 133 -77
rect 126 -80 133 -79
rect 163 -63 170 -62
rect 163 -65 165 -63
rect 167 -65 170 -63
rect 163 -66 170 -65
rect 174 -65 178 -63
rect 174 -67 175 -65
rect 177 -67 178 -65
rect 174 -77 178 -67
rect 200 -54 204 -52
rect 200 -56 201 -54
rect 203 -56 204 -54
rect 200 -60 204 -56
rect 200 -62 212 -60
rect 200 -64 207 -62
rect 209 -64 212 -62
rect 200 -66 212 -64
rect 165 -78 178 -77
rect 232 -46 236 -41
rect 232 -48 233 -46
rect 235 -48 236 -46
rect 232 -53 236 -48
rect 232 -55 233 -53
rect 235 -55 236 -53
rect 232 -76 236 -55
rect 272 -54 284 -52
rect 272 -56 280 -54
rect 282 -56 284 -54
rect 272 -58 284 -56
rect 272 -62 276 -58
rect 165 -80 167 -78
rect 169 -80 178 -78
rect 165 -81 178 -80
rect 232 -77 239 -76
rect 232 -79 235 -77
rect 237 -79 239 -77
rect 232 -80 239 -79
rect 269 -63 276 -62
rect 269 -65 271 -63
rect 273 -65 276 -63
rect 269 -66 276 -65
rect 280 -65 284 -63
rect 280 -67 281 -65
rect 283 -67 284 -65
rect 280 -77 284 -67
rect 306 -53 310 -52
rect 306 -55 307 -53
rect 309 -55 310 -53
rect 306 -60 310 -55
rect 306 -62 318 -60
rect 306 -64 313 -62
rect 315 -64 318 -62
rect 306 -66 318 -64
rect 271 -78 284 -77
rect 338 -46 342 -41
rect 338 -48 339 -46
rect 341 -48 342 -46
rect 338 -53 342 -48
rect 338 -55 339 -53
rect 341 -55 342 -53
rect 338 -76 342 -55
rect 378 -54 390 -52
rect 378 -56 386 -54
rect 388 -56 390 -54
rect 378 -58 390 -56
rect 378 -62 382 -58
rect 271 -80 273 -78
rect 275 -80 284 -78
rect 271 -81 284 -80
rect 338 -77 345 -76
rect 338 -79 341 -77
rect 343 -79 345 -77
rect 338 -80 345 -79
rect 375 -63 382 -62
rect 375 -65 377 -63
rect 379 -65 382 -63
rect 375 -66 382 -65
rect 386 -65 390 -63
rect 386 -67 387 -65
rect 389 -67 390 -65
rect 386 -77 390 -67
rect 412 -54 416 -52
rect 412 -56 413 -54
rect 415 -56 416 -54
rect 412 -60 416 -56
rect 412 -62 424 -60
rect 412 -64 419 -62
rect 421 -64 424 -62
rect 412 -66 424 -64
rect 377 -78 390 -77
rect 444 -46 448 -41
rect 444 -48 445 -46
rect 447 -48 448 -46
rect 444 -53 448 -48
rect 444 -55 445 -53
rect 447 -55 448 -53
rect 444 -76 448 -55
rect 484 -55 496 -52
rect 484 -57 491 -55
rect 493 -57 496 -55
rect 484 -58 496 -57
rect 484 -62 488 -58
rect 377 -80 379 -78
rect 381 -80 390 -78
rect 377 -81 390 -80
rect 444 -77 451 -76
rect 444 -79 447 -77
rect 449 -79 451 -77
rect 444 -80 451 -79
rect 481 -63 488 -62
rect 481 -65 483 -63
rect 485 -65 488 -63
rect 481 -66 488 -65
rect 492 -65 496 -63
rect 492 -67 493 -65
rect 495 -67 496 -65
rect 492 -77 496 -67
rect 518 -54 522 -52
rect 518 -56 519 -54
rect 521 -56 522 -54
rect 518 -60 522 -56
rect 518 -62 530 -60
rect 518 -64 525 -62
rect 527 -64 530 -62
rect 518 -66 530 -64
rect 483 -78 496 -77
rect 550 -46 554 -41
rect 550 -48 551 -46
rect 553 -48 554 -46
rect 550 -53 554 -48
rect 550 -55 551 -53
rect 553 -55 554 -53
rect 550 -76 554 -55
rect 590 -54 602 -52
rect 590 -56 598 -54
rect 600 -56 602 -54
rect 590 -58 602 -56
rect 590 -62 594 -58
rect 483 -80 485 -78
rect 487 -80 496 -78
rect 483 -81 496 -80
rect 550 -77 557 -76
rect 550 -79 553 -77
rect 555 -79 557 -77
rect 550 -80 557 -79
rect 587 -63 594 -62
rect 587 -65 589 -63
rect 591 -65 594 -63
rect 587 -66 594 -65
rect 598 -65 602 -63
rect 598 -67 599 -65
rect 601 -67 602 -65
rect 598 -77 602 -67
rect 624 -54 628 -52
rect 624 -56 625 -54
rect 627 -56 628 -54
rect 624 -60 628 -56
rect 624 -62 636 -60
rect 624 -64 631 -62
rect 633 -64 636 -62
rect 624 -66 636 -64
rect 589 -78 602 -77
rect 656 -46 660 -41
rect 656 -48 657 -46
rect 659 -48 660 -46
rect 656 -53 660 -48
rect 656 -55 657 -53
rect 659 -55 660 -53
rect 656 -76 660 -55
rect 696 -54 708 -52
rect 696 -56 702 -54
rect 704 -56 708 -54
rect 696 -58 708 -56
rect 696 -62 700 -58
rect 589 -80 591 -78
rect 593 -80 602 -78
rect 589 -81 602 -80
rect 656 -77 663 -76
rect 656 -79 659 -77
rect 661 -79 663 -77
rect 656 -80 663 -79
rect 693 -63 700 -62
rect 693 -65 695 -63
rect 697 -65 700 -63
rect 693 -66 700 -65
rect 704 -65 708 -63
rect 704 -67 705 -65
rect 707 -67 708 -65
rect 704 -77 708 -67
rect 730 -55 734 -52
rect 730 -57 731 -55
rect 733 -57 734 -55
rect 730 -60 734 -57
rect 730 -62 742 -60
rect 730 -64 737 -62
rect 739 -64 742 -62
rect 730 -66 742 -64
rect 695 -78 708 -77
rect 762 -46 766 -41
rect 762 -48 763 -46
rect 765 -48 766 -46
rect 762 -53 766 -48
rect 762 -55 763 -53
rect 765 -55 766 -53
rect 762 -76 766 -55
rect 802 -54 814 -52
rect 802 -56 809 -54
rect 811 -56 814 -54
rect 802 -58 814 -56
rect 802 -62 806 -58
rect 695 -80 697 -78
rect 699 -80 708 -78
rect 695 -81 708 -80
rect 762 -77 769 -76
rect 762 -79 765 -77
rect 767 -79 769 -77
rect 762 -80 769 -79
rect 799 -63 806 -62
rect 799 -65 801 -63
rect 803 -65 806 -63
rect 799 -66 806 -65
rect 810 -65 814 -63
rect 810 -67 811 -65
rect 813 -67 814 -65
rect 810 -77 814 -67
rect 801 -78 814 -77
rect 827 -56 840 -52
rect 801 -80 803 -78
rect 805 -80 814 -78
rect 801 -81 814 -80
rect 827 -87 832 -56
rect 836 -60 840 -56
rect 836 -62 848 -60
rect 836 -64 843 -62
rect 845 -64 848 -62
rect 836 -66 848 -64
rect 868 -46 872 -41
rect 868 -48 869 -46
rect 871 -48 872 -46
rect 868 -53 872 -48
rect 868 -55 869 -53
rect 871 -55 872 -53
rect 868 -76 872 -55
rect 908 -54 920 -52
rect 908 -56 916 -54
rect 918 -56 920 -54
rect 908 -58 920 -56
rect 908 -62 912 -58
rect 868 -77 875 -76
rect 868 -79 871 -77
rect 873 -79 875 -77
rect 868 -80 875 -79
rect 905 -63 912 -62
rect 905 -65 907 -63
rect 909 -65 912 -63
rect 905 -66 912 -65
rect 916 -65 920 -63
rect 916 -67 917 -65
rect 919 -67 920 -65
rect 916 -77 920 -67
rect 907 -78 920 -77
rect 907 -80 909 -78
rect 911 -80 920 -78
rect 907 -81 920 -80
rect -16 -88 932 -87
rect -16 -90 -9 -88
rect -7 -90 -2 -88
rect 0 -90 97 -88
rect 99 -90 104 -88
rect 106 -90 203 -88
rect 205 -90 210 -88
rect 212 -90 309 -88
rect 311 -90 316 -88
rect 318 -90 415 -88
rect 417 -90 422 -88
rect 424 -90 521 -88
rect 523 -90 528 -88
rect 530 -90 627 -88
rect 629 -90 634 -88
rect 636 -90 733 -88
rect 735 -90 740 -88
rect 742 -90 839 -88
rect 841 -90 846 -88
rect 848 -90 932 -88
rect -16 -95 932 -90
<< alu2 >>
rect 298 1174 377 1175
rect 192 1172 240 1173
rect 192 1170 193 1172
rect 195 1170 240 1172
rect 298 1172 299 1174
rect 301 1172 377 1174
rect 298 1171 377 1172
rect 192 1169 240 1170
rect 88 1165 92 1167
rect 88 1163 89 1165
rect 91 1163 92 1165
rect 136 1166 168 1167
rect 136 1164 137 1166
rect 139 1164 165 1166
rect 167 1164 168 1166
rect 236 1166 240 1169
rect 236 1164 237 1166
rect 239 1164 240 1166
rect 314 1166 326 1167
rect 136 1163 168 1164
rect 209 1163 213 1164
rect 236 1163 240 1164
rect 284 1163 288 1165
rect 314 1164 315 1166
rect 317 1164 323 1166
rect 325 1164 326 1166
rect 314 1163 326 1164
rect 338 1163 351 1164
rect 50 1142 84 1143
rect 50 1140 81 1142
rect 83 1140 84 1142
rect 50 1139 84 1140
rect 50 1013 54 1139
rect 80 1070 84 1071
rect 80 1068 81 1070
rect 83 1068 84 1070
rect 80 1055 84 1068
rect 80 1053 81 1055
rect 83 1053 84 1055
rect 80 1052 84 1053
rect 50 1011 51 1013
rect 53 1011 54 1013
rect 50 1004 54 1011
rect 88 1021 92 1163
rect 209 1161 210 1163
rect 212 1161 213 1163
rect 209 1159 213 1161
rect 284 1161 285 1163
rect 287 1161 288 1163
rect 338 1161 339 1163
rect 341 1161 348 1163
rect 350 1161 351 1163
rect 284 1159 288 1161
rect 306 1160 310 1161
rect 338 1160 351 1161
rect 209 1157 210 1159
rect 212 1157 213 1159
rect 209 1156 213 1157
rect 306 1158 307 1160
rect 309 1158 310 1160
rect 88 1019 89 1021
rect 91 1019 92 1021
rect 31 998 84 999
rect 31 996 81 998
rect 83 996 84 998
rect 31 995 84 996
rect 31 719 35 995
rect 50 985 54 987
rect 50 983 51 985
rect 53 983 54 985
rect 50 722 54 983
rect 80 928 84 929
rect 80 926 81 928
rect 83 926 84 928
rect 80 924 84 926
rect 80 922 81 924
rect 83 922 84 924
rect 80 921 84 922
rect 77 916 81 917
rect 77 914 78 916
rect 80 914 81 916
rect 77 878 81 914
rect 77 876 78 878
rect 80 876 81 878
rect 77 875 81 876
rect 50 720 51 722
rect 53 720 54 722
rect 50 719 54 720
rect 88 733 92 1019
rect 96 1149 168 1150
rect 96 1147 165 1149
rect 167 1147 168 1149
rect 96 1146 168 1147
rect 96 1068 100 1146
rect 104 1141 136 1142
rect 306 1141 310 1158
rect 373 1158 377 1171
rect 683 1173 733 1174
rect 683 1171 730 1173
rect 732 1171 733 1173
rect 683 1170 733 1171
rect 683 1166 687 1170
rect 683 1164 684 1166
rect 686 1164 687 1166
rect 660 1162 664 1164
rect 683 1163 687 1164
rect 729 1165 733 1166
rect 729 1163 730 1165
rect 732 1163 733 1165
rect 373 1156 374 1158
rect 376 1156 377 1158
rect 373 1155 377 1156
rect 547 1157 598 1161
rect 660 1160 661 1162
rect 663 1160 664 1162
rect 660 1158 664 1160
rect 338 1148 381 1149
rect 338 1146 339 1148
rect 341 1146 381 1148
rect 338 1145 381 1146
rect 104 1139 133 1141
rect 135 1139 136 1141
rect 104 1138 136 1139
rect 216 1140 220 1141
rect 216 1138 217 1140
rect 219 1138 220 1140
rect 104 1086 108 1138
rect 153 1136 157 1137
rect 153 1134 154 1136
rect 156 1134 157 1136
rect 104 1084 105 1086
rect 107 1084 108 1086
rect 104 1083 108 1084
rect 132 1130 157 1134
rect 132 1078 136 1130
rect 216 1128 220 1138
rect 306 1137 340 1141
rect 234 1132 268 1133
rect 234 1130 235 1132
rect 237 1130 268 1132
rect 234 1129 268 1130
rect 181 1124 220 1128
rect 144 1107 148 1108
rect 144 1105 145 1107
rect 147 1105 148 1107
rect 144 1091 148 1105
rect 144 1089 145 1091
rect 147 1089 148 1091
rect 144 1087 148 1089
rect 163 1085 171 1086
rect 163 1083 164 1085
rect 166 1083 168 1085
rect 170 1083 171 1085
rect 163 1082 171 1083
rect 132 1076 133 1078
rect 135 1076 136 1078
rect 132 1074 136 1076
rect 168 1071 177 1072
rect 168 1069 169 1071
rect 171 1069 174 1071
rect 176 1069 177 1071
rect 168 1068 177 1069
rect 96 1066 97 1068
rect 99 1066 100 1068
rect 96 865 100 1066
rect 181 1061 185 1124
rect 201 1107 260 1108
rect 201 1105 202 1107
rect 204 1105 260 1107
rect 201 1104 260 1105
rect 256 1101 260 1104
rect 256 1099 257 1101
rect 259 1099 260 1101
rect 256 1098 260 1099
rect 197 1093 254 1094
rect 197 1091 198 1093
rect 200 1091 254 1093
rect 197 1090 254 1091
rect 264 1093 268 1129
rect 336 1107 340 1137
rect 336 1105 337 1107
rect 339 1105 340 1107
rect 336 1104 340 1105
rect 366 1140 370 1141
rect 366 1138 367 1140
rect 369 1138 370 1140
rect 264 1091 265 1093
rect 267 1091 268 1093
rect 264 1090 268 1091
rect 250 1086 254 1090
rect 220 1085 224 1086
rect 220 1083 221 1085
rect 223 1083 224 1085
rect 116 1060 185 1061
rect 116 1058 117 1060
rect 119 1058 185 1060
rect 116 1057 185 1058
rect 212 1068 216 1069
rect 212 1066 213 1068
rect 215 1066 216 1068
rect 156 1037 160 1057
rect 212 1047 216 1066
rect 212 1045 213 1047
rect 215 1045 216 1047
rect 212 1044 216 1045
rect 220 1047 224 1083
rect 250 1085 276 1086
rect 250 1083 273 1085
rect 275 1083 276 1085
rect 250 1082 276 1083
rect 229 1071 233 1072
rect 366 1071 370 1138
rect 229 1069 230 1071
rect 232 1069 233 1071
rect 320 1070 370 1071
rect 229 1068 233 1069
rect 229 1066 230 1068
rect 232 1066 233 1068
rect 229 1055 233 1066
rect 297 1069 301 1070
rect 297 1067 298 1069
rect 300 1067 301 1069
rect 320 1068 321 1070
rect 323 1068 370 1070
rect 320 1067 370 1068
rect 297 1063 301 1067
rect 297 1062 348 1063
rect 297 1060 345 1062
rect 347 1060 348 1062
rect 297 1059 348 1060
rect 229 1054 340 1055
rect 229 1052 337 1054
rect 339 1052 340 1054
rect 229 1051 340 1052
rect 220 1045 221 1047
rect 223 1045 224 1047
rect 220 1044 224 1045
rect 156 1035 157 1037
rect 159 1035 160 1037
rect 156 1033 160 1035
rect 203 1029 308 1030
rect 133 1028 199 1029
rect 133 1026 134 1028
rect 136 1026 199 1028
rect 203 1027 204 1029
rect 206 1027 305 1029
rect 307 1027 308 1029
rect 203 1026 308 1027
rect 133 1025 199 1026
rect 195 1021 199 1025
rect 377 1022 381 1145
rect 104 1020 164 1021
rect 104 1018 137 1020
rect 139 1018 161 1020
rect 163 1018 164 1020
rect 195 1019 196 1021
rect 198 1019 199 1021
rect 195 1018 199 1019
rect 272 1021 381 1022
rect 272 1019 273 1021
rect 275 1019 381 1021
rect 272 1018 381 1019
rect 104 1017 164 1018
rect 104 942 108 1017
rect 289 1013 373 1014
rect 289 1011 290 1013
rect 292 1011 370 1013
rect 372 1011 373 1013
rect 289 1010 373 1011
rect 236 1005 260 1006
rect 104 940 105 942
rect 107 940 108 942
rect 104 939 108 940
rect 140 1004 171 1005
rect 140 1002 168 1004
rect 170 1002 171 1004
rect 236 1003 237 1005
rect 239 1003 260 1005
rect 236 1002 260 1003
rect 140 1001 171 1002
rect 140 935 144 1001
rect 244 997 252 998
rect 148 996 152 997
rect 148 994 149 996
rect 151 994 152 996
rect 244 995 245 997
rect 247 995 252 997
rect 244 994 252 995
rect 148 963 152 994
rect 148 961 149 963
rect 151 961 152 963
rect 148 960 152 961
rect 248 957 252 994
rect 256 964 260 1002
rect 271 997 275 998
rect 271 995 272 997
rect 274 995 275 997
rect 271 993 275 995
rect 271 991 272 993
rect 274 991 275 993
rect 271 990 275 991
rect 256 960 303 964
rect 248 955 249 957
rect 251 955 252 957
rect 248 953 252 955
rect 268 950 275 951
rect 148 949 180 950
rect 148 947 149 949
rect 151 947 177 949
rect 179 947 180 949
rect 268 948 269 950
rect 271 948 272 950
rect 274 948 275 950
rect 268 947 275 948
rect 148 946 180 947
rect 299 946 303 960
rect 308 950 364 951
rect 308 948 309 950
rect 311 948 364 950
rect 308 947 364 948
rect 299 944 300 946
rect 302 944 303 946
rect 299 943 303 944
rect 104 934 144 935
rect 104 932 105 934
rect 107 932 144 934
rect 104 931 144 932
rect 200 934 204 937
rect 200 932 201 934
rect 203 932 204 934
rect 200 931 204 932
rect 144 925 243 926
rect 104 924 128 925
rect 104 922 105 924
rect 107 922 121 924
rect 123 922 125 924
rect 127 922 128 924
rect 144 923 145 925
rect 147 923 240 925
rect 242 923 243 925
rect 144 922 243 923
rect 269 924 280 925
rect 269 922 270 924
rect 272 922 277 924
rect 279 922 280 924
rect 104 921 128 922
rect 269 921 280 922
rect 116 916 189 917
rect 116 914 117 916
rect 119 914 185 916
rect 187 914 189 916
rect 116 913 189 914
rect 120 901 348 902
rect 120 899 121 901
rect 123 899 345 901
rect 347 899 348 901
rect 120 898 348 899
rect 148 891 328 892
rect 148 889 149 891
rect 151 889 325 891
rect 327 889 328 891
rect 148 888 328 889
rect 156 883 160 884
rect 156 881 157 883
rect 159 881 160 883
rect 105 878 145 879
rect 105 876 106 878
rect 108 876 141 878
rect 143 876 145 878
rect 105 875 145 876
rect 96 863 97 865
rect 99 863 100 865
rect 96 862 100 863
rect 139 861 143 862
rect 139 859 140 861
rect 142 859 143 861
rect 139 857 143 859
rect 101 853 143 857
rect 101 809 105 853
rect 116 847 143 848
rect 116 845 117 847
rect 119 845 143 847
rect 116 844 143 845
rect 101 807 102 809
rect 104 807 105 809
rect 101 806 105 807
rect 112 839 116 840
rect 112 837 113 839
rect 115 837 116 839
rect 112 806 116 837
rect 112 804 113 806
rect 115 804 116 806
rect 112 803 116 804
rect 116 797 120 798
rect 116 795 117 797
rect 119 795 120 797
rect 88 731 89 733
rect 91 731 92 733
rect 31 717 32 719
rect 34 717 35 719
rect 31 716 35 717
rect 20 711 84 712
rect 20 709 81 711
rect 83 709 84 711
rect 20 708 84 709
rect 20 582 24 708
rect 50 703 54 704
rect 50 701 51 703
rect 53 701 54 703
rect 31 692 35 694
rect 31 690 32 692
rect 34 690 35 692
rect 31 589 35 690
rect 31 587 32 589
rect 34 587 35 589
rect 31 582 35 587
rect 20 580 21 582
rect 23 580 24 582
rect 20 578 24 580
rect 50 581 54 701
rect 88 608 92 731
rect 96 781 100 782
rect 96 779 97 781
rect 99 779 100 781
rect 96 777 100 779
rect 96 775 97 777
rect 99 775 100 777
rect 96 658 100 775
rect 116 772 120 795
rect 139 789 143 844
rect 156 804 160 881
rect 180 883 320 884
rect 180 881 181 883
rect 183 881 320 883
rect 180 880 320 881
rect 316 878 320 880
rect 316 876 317 878
rect 319 876 320 878
rect 189 875 224 876
rect 189 873 190 875
rect 192 873 221 875
rect 223 873 224 875
rect 189 872 224 873
rect 254 875 268 876
rect 316 875 320 876
rect 254 873 255 875
rect 257 873 265 875
rect 267 873 268 875
rect 254 872 268 873
rect 228 869 232 870
rect 228 867 229 869
rect 231 867 232 869
rect 156 802 157 804
rect 159 802 160 804
rect 156 801 160 802
rect 165 856 169 857
rect 165 854 166 856
rect 168 854 169 856
rect 139 787 140 789
rect 142 787 143 789
rect 139 786 143 787
rect 165 785 169 854
rect 211 853 222 854
rect 197 852 207 853
rect 197 850 198 852
rect 200 850 204 852
rect 206 850 207 852
rect 197 849 207 850
rect 211 851 219 853
rect 221 851 222 853
rect 211 850 222 851
rect 180 839 184 840
rect 180 837 181 839
rect 183 837 184 839
rect 180 806 184 837
rect 180 804 181 806
rect 183 804 184 806
rect 180 803 184 804
rect 197 819 201 820
rect 197 817 198 819
rect 200 817 201 819
rect 197 789 201 817
rect 211 803 215 850
rect 211 801 212 803
rect 214 801 215 803
rect 211 800 215 801
rect 228 803 232 867
rect 280 868 284 869
rect 280 866 281 868
rect 283 866 284 868
rect 280 865 284 866
rect 250 864 284 865
rect 250 862 251 864
rect 253 862 284 864
rect 250 861 284 862
rect 324 861 328 888
rect 324 859 325 861
rect 327 859 328 861
rect 324 858 328 859
rect 360 869 364 947
rect 360 867 361 869
rect 363 867 364 869
rect 292 856 296 857
rect 292 854 293 856
rect 295 854 296 856
rect 292 840 296 854
rect 337 845 341 846
rect 337 843 338 845
rect 340 843 341 845
rect 228 801 229 803
rect 231 801 232 803
rect 228 800 232 801
rect 269 839 273 840
rect 269 837 270 839
rect 272 837 273 839
rect 269 799 273 837
rect 292 836 320 840
rect 280 819 284 820
rect 280 817 281 819
rect 283 817 284 819
rect 280 806 284 817
rect 280 804 281 806
rect 283 804 284 806
rect 280 803 284 804
rect 260 798 279 799
rect 260 796 261 798
rect 263 796 276 798
rect 278 796 279 798
rect 260 795 279 796
rect 197 787 198 789
rect 200 787 201 789
rect 197 786 201 787
rect 316 789 320 836
rect 337 807 341 843
rect 333 806 341 807
rect 333 804 334 806
rect 336 804 341 806
rect 333 803 341 804
rect 316 787 317 789
rect 319 787 320 789
rect 316 786 320 787
rect 165 783 166 785
rect 168 783 169 785
rect 165 781 169 783
rect 253 780 257 781
rect 253 778 254 780
rect 256 778 257 780
rect 116 770 117 772
rect 119 770 120 772
rect 116 769 120 770
rect 124 772 128 773
rect 124 770 125 772
rect 127 770 128 772
rect 124 747 128 770
rect 253 768 257 778
rect 280 780 305 781
rect 280 778 281 780
rect 283 778 302 780
rect 304 778 305 780
rect 280 777 305 778
rect 360 768 364 867
rect 124 745 125 747
rect 127 745 128 747
rect 124 744 128 745
rect 215 764 364 768
rect 369 853 373 1010
rect 369 851 370 853
rect 372 851 373 853
rect 136 741 197 742
rect 136 739 137 741
rect 139 739 197 741
rect 136 738 197 739
rect 193 725 197 738
rect 148 724 152 725
rect 148 722 149 724
rect 151 722 152 724
rect 193 723 194 725
rect 196 723 197 725
rect 193 722 197 723
rect 215 725 219 764
rect 262 747 332 748
rect 262 745 263 747
rect 265 745 332 747
rect 262 744 332 745
rect 240 733 266 734
rect 328 733 332 744
rect 240 731 241 733
rect 243 731 263 733
rect 265 731 266 733
rect 240 730 266 731
rect 308 731 312 733
rect 308 729 309 731
rect 311 729 312 731
rect 328 731 329 733
rect 331 731 332 733
rect 328 730 332 731
rect 308 727 312 729
rect 215 723 216 725
rect 218 723 219 725
rect 96 656 97 658
rect 99 656 100 658
rect 96 630 100 656
rect 113 709 135 710
rect 113 707 132 709
rect 134 707 135 709
rect 113 706 135 707
rect 113 654 117 706
rect 148 702 152 722
rect 215 718 219 723
rect 176 717 219 718
rect 176 715 177 717
rect 179 715 219 717
rect 176 714 219 715
rect 113 652 114 654
rect 116 652 117 654
rect 113 651 117 652
rect 124 698 152 702
rect 208 709 212 710
rect 208 707 209 709
rect 211 707 212 709
rect 124 638 128 698
rect 208 676 212 707
rect 328 709 365 711
rect 328 707 329 709
rect 331 707 365 709
rect 328 706 365 707
rect 146 672 212 676
rect 253 700 257 701
rect 253 698 254 700
rect 256 698 257 700
rect 146 657 150 672
rect 157 661 218 662
rect 157 659 158 661
rect 160 659 218 661
rect 253 660 257 698
rect 157 658 218 659
rect 146 655 147 657
rect 149 655 150 657
rect 146 654 150 655
rect 192 653 196 654
rect 192 651 193 653
rect 195 651 196 653
rect 105 637 128 638
rect 105 635 106 637
rect 108 635 128 637
rect 105 634 128 635
rect 132 645 136 646
rect 132 643 133 645
rect 135 643 136 645
rect 132 630 136 643
rect 96 626 136 630
rect 184 637 188 638
rect 184 635 185 637
rect 187 635 188 637
rect 184 623 188 635
rect 184 621 185 623
rect 187 621 188 623
rect 184 620 188 621
rect 192 624 196 651
rect 214 637 218 658
rect 222 659 257 660
rect 222 657 223 659
rect 225 657 257 659
rect 222 656 257 657
rect 275 683 279 684
rect 275 681 276 683
rect 278 681 279 683
rect 275 646 279 681
rect 214 635 215 637
rect 217 635 218 637
rect 214 634 218 635
rect 264 645 279 646
rect 264 643 265 645
rect 267 643 279 645
rect 264 642 279 643
rect 192 623 250 624
rect 192 621 247 623
rect 249 621 250 623
rect 192 620 250 621
rect 88 607 260 608
rect 88 605 257 607
rect 259 605 260 607
rect 88 604 260 605
rect 88 590 92 604
rect 148 598 197 599
rect 148 596 149 598
rect 151 596 185 598
rect 187 596 197 598
rect 148 595 197 596
rect 193 590 197 595
rect 88 588 89 590
rect 91 588 92 590
rect 88 587 92 588
rect 136 589 160 590
rect 136 587 137 589
rect 139 587 157 589
rect 159 587 160 589
rect 193 588 194 590
rect 196 588 197 590
rect 193 587 197 588
rect 136 586 160 587
rect 50 579 51 581
rect 53 579 54 581
rect 50 574 54 579
rect 246 582 250 583
rect 246 580 247 582
rect 249 580 250 582
rect 246 577 250 580
rect 199 575 222 576
rect 199 573 219 575
rect 221 573 222 575
rect 165 572 169 573
rect 165 570 166 572
rect 168 570 169 572
rect 5 567 84 568
rect 5 565 81 567
rect 83 565 84 567
rect 5 564 84 565
rect 90 564 133 565
rect 5 335 9 564
rect 90 562 130 564
rect 132 562 133 564
rect 90 561 133 562
rect 20 554 24 558
rect 20 552 21 554
rect 23 552 24 554
rect 20 379 24 552
rect 31 552 35 554
rect 31 550 32 552
rect 34 550 35 552
rect 31 389 35 550
rect 50 553 54 555
rect 50 551 51 553
rect 53 551 54 553
rect 50 398 54 551
rect 80 551 84 552
rect 80 549 81 551
rect 83 549 84 551
rect 80 509 84 549
rect 80 507 81 509
rect 83 507 84 509
rect 80 506 84 507
rect 90 493 94 561
rect 165 557 169 570
rect 199 572 222 573
rect 246 575 247 577
rect 249 575 250 577
rect 113 553 169 557
rect 186 564 190 565
rect 186 562 187 564
rect 189 562 190 564
rect 113 510 117 553
rect 186 517 190 562
rect 138 516 190 517
rect 138 514 139 516
rect 141 514 190 516
rect 138 513 190 514
rect 113 508 114 510
rect 116 508 117 510
rect 113 507 117 508
rect 199 502 203 572
rect 238 565 242 567
rect 238 563 239 565
rect 241 563 242 565
rect 238 527 242 563
rect 215 526 242 527
rect 215 524 216 526
rect 218 524 242 526
rect 215 523 242 524
rect 246 517 250 575
rect 246 515 247 517
rect 249 515 250 517
rect 246 514 250 515
rect 256 510 260 604
rect 264 551 268 642
rect 361 616 365 706
rect 369 632 373 851
rect 369 630 370 632
rect 372 630 373 632
rect 369 629 373 630
rect 377 878 381 1018
rect 377 876 378 878
rect 380 876 381 878
rect 377 623 381 876
rect 377 621 378 623
rect 380 621 381 623
rect 377 620 381 621
rect 400 1040 507 1044
rect 400 616 404 1040
rect 361 612 404 616
rect 389 611 404 612
rect 442 1035 446 1036
rect 442 1033 443 1035
rect 445 1033 446 1035
rect 442 780 446 1033
rect 442 778 443 780
rect 445 778 446 780
rect 442 638 446 778
rect 450 1026 454 1027
rect 450 1024 451 1026
rect 453 1024 454 1026
rect 450 805 454 1024
rect 503 1015 507 1040
rect 547 1031 551 1157
rect 594 1150 598 1157
rect 590 1149 598 1150
rect 590 1147 591 1149
rect 593 1147 598 1149
rect 590 1146 598 1147
rect 620 1156 624 1157
rect 620 1154 621 1156
rect 623 1154 624 1156
rect 573 1141 577 1142
rect 573 1139 574 1141
rect 576 1139 577 1141
rect 511 1030 551 1031
rect 511 1028 512 1030
rect 514 1028 551 1030
rect 511 1027 551 1028
rect 555 1107 559 1108
rect 555 1105 556 1107
rect 558 1105 559 1107
rect 503 1014 531 1015
rect 555 1014 559 1105
rect 573 1081 577 1139
rect 581 1132 608 1133
rect 581 1130 605 1132
rect 607 1130 608 1132
rect 581 1129 608 1130
rect 581 1093 585 1129
rect 581 1091 582 1093
rect 584 1091 585 1093
rect 581 1089 585 1091
rect 620 1084 624 1154
rect 706 1148 710 1149
rect 706 1146 707 1148
rect 709 1146 710 1148
rect 633 1142 685 1143
rect 633 1140 682 1142
rect 684 1140 685 1142
rect 633 1139 685 1140
rect 633 1094 637 1139
rect 706 1103 710 1146
rect 633 1092 634 1094
rect 636 1092 637 1094
rect 633 1091 637 1092
rect 654 1099 710 1103
rect 573 1079 574 1081
rect 576 1079 577 1081
rect 601 1083 624 1084
rect 654 1086 658 1099
rect 729 1095 733 1163
rect 739 1149 743 1150
rect 739 1147 740 1149
rect 742 1147 743 1149
rect 739 1107 743 1147
rect 739 1105 740 1107
rect 742 1105 743 1107
rect 739 1104 743 1105
rect 690 1094 733 1095
rect 690 1092 691 1094
rect 693 1092 733 1094
rect 690 1091 733 1092
rect 739 1093 770 1094
rect 739 1091 740 1093
rect 742 1091 766 1093
rect 768 1091 770 1093
rect 739 1090 770 1091
rect 654 1084 655 1086
rect 657 1084 658 1086
rect 654 1083 658 1084
rect 601 1081 602 1083
rect 604 1081 624 1083
rect 601 1080 624 1081
rect 573 1076 577 1079
rect 573 1074 574 1076
rect 576 1074 577 1076
rect 573 1073 577 1074
rect 663 1069 687 1070
rect 626 1068 630 1069
rect 626 1066 627 1068
rect 629 1066 630 1068
rect 663 1067 664 1069
rect 666 1067 684 1069
rect 686 1067 687 1069
rect 663 1066 687 1067
rect 731 1068 735 1069
rect 731 1066 732 1068
rect 734 1066 735 1068
rect 626 1061 630 1066
rect 626 1060 675 1061
rect 626 1058 636 1060
rect 638 1058 672 1060
rect 674 1058 675 1060
rect 626 1057 675 1058
rect 731 1052 735 1066
rect 563 1051 735 1052
rect 563 1049 564 1051
rect 566 1049 735 1051
rect 563 1048 735 1049
rect 573 1035 631 1036
rect 573 1033 574 1035
rect 576 1033 631 1035
rect 573 1032 631 1033
rect 503 1012 528 1014
rect 530 1012 531 1014
rect 503 1011 531 1012
rect 544 1013 559 1014
rect 544 1011 556 1013
rect 558 1011 559 1013
rect 544 1010 559 1011
rect 605 1021 609 1022
rect 605 1019 606 1021
rect 608 1019 609 1021
rect 544 975 548 1010
rect 544 973 545 975
rect 547 973 548 975
rect 544 972 548 973
rect 566 999 601 1000
rect 566 997 598 999
rect 600 997 601 999
rect 566 996 601 997
rect 605 998 609 1019
rect 627 1005 631 1032
rect 635 1035 639 1036
rect 635 1033 636 1035
rect 638 1033 639 1035
rect 635 1021 639 1033
rect 635 1019 636 1021
rect 638 1019 639 1021
rect 635 1018 639 1019
rect 687 1026 727 1030
rect 687 1013 691 1026
rect 687 1011 688 1013
rect 690 1011 691 1013
rect 687 1010 691 1011
rect 695 1021 718 1022
rect 695 1019 715 1021
rect 717 1019 718 1021
rect 695 1018 718 1019
rect 627 1003 628 1005
rect 630 1003 631 1005
rect 627 1002 631 1003
rect 673 1001 677 1002
rect 673 999 674 1001
rect 676 999 677 1001
rect 605 997 666 998
rect 566 958 570 996
rect 605 995 663 997
rect 665 995 666 997
rect 605 994 666 995
rect 673 984 677 999
rect 566 956 567 958
rect 569 956 570 958
rect 566 955 570 956
rect 611 980 677 984
rect 611 949 615 980
rect 695 958 699 1018
rect 611 947 612 949
rect 614 947 615 949
rect 611 946 615 947
rect 671 954 699 958
rect 706 1004 710 1005
rect 706 1002 707 1004
rect 709 1002 710 1004
rect 604 941 647 942
rect 604 939 644 941
rect 646 939 647 941
rect 604 938 647 939
rect 604 933 608 938
rect 671 934 675 954
rect 706 950 710 1002
rect 688 949 710 950
rect 688 947 689 949
rect 691 947 710 949
rect 688 946 710 947
rect 723 1000 727 1026
rect 723 998 724 1000
rect 726 998 727 1000
rect 604 931 605 933
rect 607 931 608 933
rect 511 926 515 929
rect 511 924 512 926
rect 514 924 515 926
rect 511 922 515 924
rect 557 925 583 926
rect 557 923 558 925
rect 560 923 580 925
rect 582 923 583 925
rect 557 922 583 923
rect 604 892 608 931
rect 626 933 630 934
rect 626 931 627 933
rect 629 931 630 933
rect 671 932 672 934
rect 674 932 675 934
rect 671 931 675 932
rect 626 918 630 931
rect 626 917 687 918
rect 626 915 684 917
rect 686 915 687 917
rect 626 914 687 915
rect 450 803 451 805
rect 453 803 454 805
rect 450 646 454 803
rect 459 888 608 892
rect 459 789 463 888
rect 518 878 543 879
rect 518 876 519 878
rect 521 876 540 878
rect 542 876 543 878
rect 518 875 543 876
rect 566 878 570 888
rect 566 876 567 878
rect 569 876 570 878
rect 566 875 570 876
rect 703 886 707 887
rect 703 884 704 886
rect 706 884 707 886
rect 654 873 658 875
rect 654 871 655 873
rect 657 871 658 873
rect 503 869 507 870
rect 503 867 504 869
rect 506 867 507 869
rect 482 852 490 853
rect 482 850 487 852
rect 489 850 490 852
rect 482 849 490 850
rect 482 813 486 849
rect 503 820 507 867
rect 622 869 626 870
rect 622 867 623 869
rect 625 867 626 869
rect 544 860 563 861
rect 544 858 545 860
rect 547 858 560 860
rect 562 858 563 860
rect 544 857 563 858
rect 539 852 543 853
rect 539 850 540 852
rect 542 850 543 852
rect 539 839 543 850
rect 539 837 540 839
rect 542 837 543 839
rect 539 836 543 837
rect 503 816 531 820
rect 550 819 554 857
rect 550 817 551 819
rect 553 817 554 819
rect 550 816 554 817
rect 591 855 595 856
rect 591 853 592 855
rect 594 853 595 855
rect 482 811 483 813
rect 485 811 486 813
rect 482 810 486 811
rect 527 802 531 816
rect 527 800 528 802
rect 530 800 531 802
rect 527 799 531 800
rect 459 787 460 789
rect 462 787 463 789
rect 459 709 463 787
rect 495 797 499 798
rect 495 795 496 797
rect 498 795 499 797
rect 495 768 499 795
rect 539 794 573 795
rect 539 792 570 794
rect 572 792 573 794
rect 539 791 573 792
rect 539 790 543 791
rect 539 788 540 790
rect 542 788 543 790
rect 539 787 543 788
rect 591 789 595 853
rect 608 855 612 856
rect 608 853 609 855
rect 611 853 612 855
rect 608 806 612 853
rect 622 839 626 867
rect 622 837 623 839
rect 625 837 626 839
rect 622 836 626 837
rect 639 852 643 853
rect 639 850 640 852
rect 642 850 643 852
rect 639 819 643 850
rect 639 817 640 819
rect 642 817 643 819
rect 639 816 643 817
rect 601 805 612 806
rect 601 803 602 805
rect 604 803 612 805
rect 616 806 626 807
rect 616 804 617 806
rect 619 804 623 806
rect 625 804 626 806
rect 616 803 626 804
rect 601 802 612 803
rect 654 802 658 871
rect 680 869 684 870
rect 680 867 681 869
rect 683 867 684 869
rect 654 800 655 802
rect 657 800 658 802
rect 654 799 658 800
rect 663 854 667 855
rect 663 852 664 854
rect 666 852 667 854
rect 591 787 592 789
rect 594 787 595 789
rect 591 786 595 787
rect 555 783 569 784
rect 555 781 556 783
rect 558 781 566 783
rect 568 781 569 783
rect 503 780 507 781
rect 555 780 569 781
rect 599 783 634 784
rect 599 781 600 783
rect 602 781 631 783
rect 633 781 634 783
rect 599 780 634 781
rect 503 778 504 780
rect 506 778 507 780
rect 503 776 507 778
rect 503 775 643 776
rect 503 773 640 775
rect 642 773 643 775
rect 503 772 643 773
rect 663 775 667 852
rect 680 812 684 867
rect 695 867 699 869
rect 695 865 696 867
rect 698 865 699 867
rect 695 862 699 865
rect 703 861 707 884
rect 723 881 727 998
rect 723 879 724 881
rect 726 879 727 881
rect 723 877 727 879
rect 723 875 724 877
rect 726 875 727 877
rect 723 874 727 875
rect 731 925 735 1048
rect 739 949 816 950
rect 739 947 740 949
rect 742 947 816 949
rect 739 946 816 947
rect 731 923 732 925
rect 734 923 735 925
rect 703 859 704 861
rect 706 859 707 861
rect 703 858 707 859
rect 707 852 711 853
rect 707 850 708 852
rect 710 850 711 852
rect 707 819 711 850
rect 707 817 708 819
rect 710 817 711 819
rect 707 816 711 817
rect 718 849 722 850
rect 718 847 719 849
rect 721 847 722 849
rect 680 811 707 812
rect 680 809 704 811
rect 706 809 707 811
rect 680 808 707 809
rect 718 803 722 847
rect 680 799 722 803
rect 680 797 684 799
rect 680 795 681 797
rect 683 795 684 797
rect 680 794 684 795
rect 723 793 727 794
rect 723 791 724 793
rect 726 791 727 793
rect 678 780 718 781
rect 678 778 680 780
rect 682 778 715 780
rect 717 778 718 780
rect 678 777 718 778
rect 663 773 664 775
rect 666 773 667 775
rect 663 772 667 773
rect 495 767 675 768
rect 495 765 496 767
rect 498 765 672 767
rect 674 765 675 767
rect 495 764 675 765
rect 475 757 703 758
rect 475 755 476 757
rect 478 755 700 757
rect 702 755 703 757
rect 475 754 703 755
rect 634 742 707 743
rect 634 740 636 742
rect 638 740 704 742
rect 706 740 707 742
rect 634 739 707 740
rect 543 734 554 735
rect 695 734 719 735
rect 543 732 544 734
rect 546 732 551 734
rect 553 732 554 734
rect 543 731 554 732
rect 580 733 679 734
rect 580 731 581 733
rect 583 731 676 733
rect 678 731 679 733
rect 695 732 696 734
rect 698 732 700 734
rect 702 732 716 734
rect 718 732 719 734
rect 695 731 719 732
rect 580 730 679 731
rect 619 723 623 726
rect 619 721 620 723
rect 622 721 623 723
rect 619 719 623 721
rect 679 724 719 725
rect 679 722 716 724
rect 718 722 719 724
rect 679 721 719 722
rect 520 712 524 713
rect 520 710 521 712
rect 523 710 524 712
rect 459 708 515 709
rect 459 706 512 708
rect 514 706 515 708
rect 459 705 515 706
rect 520 696 524 710
rect 643 709 675 710
rect 548 708 555 709
rect 548 706 549 708
rect 551 706 552 708
rect 554 706 555 708
rect 643 707 644 709
rect 646 707 672 709
rect 674 707 675 709
rect 643 706 675 707
rect 548 705 555 706
rect 571 701 575 703
rect 571 699 572 701
rect 574 699 575 701
rect 520 692 567 696
rect 548 665 552 666
rect 548 663 549 665
rect 551 663 552 665
rect 548 661 552 663
rect 548 659 549 661
rect 551 659 552 661
rect 548 658 552 659
rect 563 654 567 692
rect 571 662 575 699
rect 671 695 675 696
rect 671 693 672 695
rect 674 693 675 695
rect 671 662 675 693
rect 571 661 579 662
rect 571 659 576 661
rect 578 659 579 661
rect 671 660 672 662
rect 674 660 675 662
rect 671 659 675 660
rect 571 658 579 659
rect 679 655 683 721
rect 652 654 683 655
rect 563 653 587 654
rect 563 651 584 653
rect 586 651 587 653
rect 652 652 653 654
rect 655 652 683 654
rect 652 651 683 652
rect 715 716 719 717
rect 715 714 716 716
rect 718 714 719 716
rect 563 650 587 651
rect 450 645 534 646
rect 450 643 451 645
rect 453 643 531 645
rect 533 643 534 645
rect 450 642 534 643
rect 715 639 719 714
rect 659 638 719 639
rect 442 637 551 638
rect 442 635 548 637
rect 550 635 551 637
rect 442 634 551 635
rect 624 637 628 638
rect 624 635 625 637
rect 627 635 628 637
rect 659 636 660 638
rect 662 636 684 638
rect 686 636 719 638
rect 659 635 719 636
rect 264 549 265 551
rect 267 549 268 551
rect 264 548 268 549
rect 238 509 260 510
rect 238 507 239 509
rect 241 507 260 509
rect 442 511 446 634
rect 624 631 628 635
rect 624 630 690 631
rect 515 629 620 630
rect 515 627 516 629
rect 518 627 617 629
rect 619 627 620 629
rect 624 628 687 630
rect 689 628 690 630
rect 624 627 690 628
rect 515 626 620 627
rect 663 621 667 623
rect 663 619 664 621
rect 666 619 667 621
rect 599 611 603 612
rect 599 609 600 611
rect 602 609 603 611
rect 483 604 594 605
rect 483 602 484 604
rect 486 602 594 604
rect 483 601 594 602
rect 475 596 526 597
rect 475 594 476 596
rect 478 594 526 596
rect 475 593 526 594
rect 522 589 526 593
rect 453 588 503 589
rect 453 586 500 588
rect 502 586 503 588
rect 522 587 523 589
rect 525 587 526 589
rect 522 586 526 587
rect 590 590 594 601
rect 590 588 591 590
rect 593 588 594 590
rect 590 587 594 588
rect 453 585 503 586
rect 590 585 591 587
rect 593 585 594 587
rect 453 518 457 585
rect 590 584 594 585
rect 547 573 573 574
rect 547 571 548 573
rect 550 571 573 573
rect 547 570 573 571
rect 599 573 603 609
rect 607 611 611 612
rect 607 609 608 611
rect 610 609 611 611
rect 607 590 611 609
rect 663 599 667 619
rect 607 588 608 590
rect 610 588 611 590
rect 607 587 611 588
rect 638 598 707 599
rect 638 596 704 598
rect 706 596 707 598
rect 638 595 707 596
rect 599 571 600 573
rect 602 571 603 573
rect 599 570 603 571
rect 569 566 573 570
rect 555 565 559 566
rect 555 563 556 565
rect 558 563 559 565
rect 453 516 454 518
rect 456 516 457 518
rect 453 515 457 516
rect 483 551 487 552
rect 483 549 484 551
rect 486 549 487 551
rect 483 519 487 549
rect 555 527 559 563
rect 569 565 626 566
rect 569 563 623 565
rect 625 563 626 565
rect 569 562 626 563
rect 563 557 567 558
rect 563 555 564 557
rect 566 555 567 557
rect 563 552 567 555
rect 563 551 622 552
rect 563 549 619 551
rect 621 549 622 551
rect 563 548 622 549
rect 638 532 642 595
rect 723 590 727 791
rect 723 588 724 590
rect 726 588 727 590
rect 646 587 655 588
rect 646 585 647 587
rect 649 585 652 587
rect 654 585 655 587
rect 646 584 655 585
rect 687 580 691 582
rect 687 578 688 580
rect 690 578 691 580
rect 652 573 660 574
rect 652 571 653 573
rect 655 571 657 573
rect 659 571 660 573
rect 652 570 660 571
rect 675 567 679 569
rect 675 565 676 567
rect 678 565 679 567
rect 675 551 679 565
rect 675 549 676 551
rect 678 549 679 551
rect 675 548 679 549
rect 603 528 642 532
rect 555 526 589 527
rect 555 524 586 526
rect 588 524 589 526
rect 555 523 589 524
rect 483 515 517 519
rect 603 518 607 528
rect 687 526 691 578
rect 666 522 691 526
rect 715 572 719 573
rect 715 570 716 572
rect 718 570 719 572
rect 666 520 667 522
rect 669 520 670 522
rect 666 519 670 520
rect 715 518 719 570
rect 603 516 604 518
rect 606 516 607 518
rect 603 515 607 516
rect 687 517 719 518
rect 687 515 688 517
rect 690 515 719 517
rect 442 510 485 511
rect 442 508 482 510
rect 484 508 485 510
rect 442 507 485 508
rect 238 506 260 507
rect 199 500 200 502
rect 202 500 203 502
rect 199 499 203 500
rect 446 500 450 501
rect 159 497 163 499
rect 159 495 160 497
rect 162 495 163 497
rect 159 493 163 495
rect 446 498 447 500
rect 449 498 450 500
rect 90 491 91 493
rect 93 491 94 493
rect 90 490 94 491
rect 136 492 140 493
rect 136 490 137 492
rect 139 490 140 492
rect 136 486 140 490
rect 90 485 140 486
rect 90 483 91 485
rect 93 483 140 485
rect 90 482 140 483
rect 446 485 450 498
rect 513 498 517 515
rect 687 514 719 515
rect 723 510 727 588
rect 655 509 727 510
rect 655 507 656 509
rect 658 507 727 509
rect 655 506 727 507
rect 731 637 735 923
rect 742 780 746 781
rect 742 778 743 780
rect 745 778 746 780
rect 742 742 746 778
rect 742 740 743 742
rect 745 740 746 742
rect 742 739 746 740
rect 739 734 743 735
rect 739 732 740 734
rect 742 732 743 734
rect 739 730 743 732
rect 739 728 740 730
rect 742 728 743 730
rect 739 727 743 728
rect 739 662 781 663
rect 739 660 740 662
rect 742 660 781 662
rect 739 659 781 660
rect 731 635 732 637
rect 734 635 735 637
rect 513 496 514 498
rect 516 496 517 498
rect 610 499 614 500
rect 610 497 611 499
rect 613 497 614 499
rect 472 495 485 496
rect 513 495 517 496
rect 535 495 539 497
rect 472 493 473 495
rect 475 493 482 495
rect 484 493 485 495
rect 535 493 536 495
rect 538 493 539 495
rect 610 495 614 497
rect 610 493 611 495
rect 613 493 614 495
rect 731 493 735 635
rect 739 603 743 604
rect 739 601 740 603
rect 742 601 743 603
rect 739 588 743 601
rect 739 586 740 588
rect 742 586 743 588
rect 739 585 743 586
rect 739 516 758 517
rect 739 514 740 516
rect 742 514 758 516
rect 739 513 758 514
rect 472 492 485 493
rect 497 492 509 493
rect 497 490 498 492
rect 500 490 506 492
rect 508 490 509 492
rect 535 491 539 493
rect 583 492 587 493
rect 610 492 614 493
rect 655 492 687 493
rect 497 489 509 490
rect 583 490 584 492
rect 586 490 587 492
rect 583 487 587 490
rect 655 490 656 492
rect 658 490 684 492
rect 686 490 687 492
rect 655 489 687 490
rect 731 491 732 493
rect 734 491 735 493
rect 731 489 735 491
rect 583 486 631 487
rect 446 484 525 485
rect 446 482 522 484
rect 524 482 525 484
rect 583 484 628 486
rect 630 484 631 486
rect 583 483 631 484
rect 446 481 525 482
rect 754 458 758 513
rect 705 457 758 458
rect 705 455 706 457
rect 708 455 758 457
rect 705 454 758 455
rect 777 436 781 659
rect 627 435 781 436
rect 627 433 630 435
rect 632 433 781 435
rect 627 432 781 433
rect 812 423 816 946
rect 500 422 816 423
rect 500 420 501 422
rect 503 420 816 422
rect 500 419 816 420
rect 50 394 125 398
rect 31 385 114 389
rect 20 378 103 379
rect 20 376 100 378
rect 102 376 103 378
rect 20 375 103 376
rect 110 375 114 385
rect 121 383 125 394
rect 121 382 271 383
rect 121 380 267 382
rect 269 380 271 382
rect 121 379 271 380
rect 110 374 205 375
rect 110 372 202 374
rect 204 372 205 374
rect 110 371 205 372
rect 77 362 705 366
rect 77 342 81 362
rect 177 354 604 358
rect 177 350 181 354
rect 600 350 604 354
rect 177 348 178 350
rect 180 348 181 350
rect 177 347 181 348
rect 201 349 205 350
rect 201 347 202 349
rect 204 347 205 349
rect 201 346 205 347
rect 277 349 504 350
rect 277 347 278 349
rect 280 347 501 349
rect 503 347 504 349
rect 600 348 601 350
rect 603 348 604 350
rect 600 347 604 348
rect 701 349 705 362
rect 701 347 702 349
rect 704 347 705 349
rect 277 346 504 347
rect 701 346 705 347
rect 77 340 78 342
rect 80 340 81 342
rect 77 339 81 340
rect 85 341 822 342
rect 85 339 86 341
rect 88 339 186 341
rect 188 339 286 341
rect 288 339 386 341
rect 388 339 486 341
rect 488 339 586 341
rect 588 339 686 341
rect 688 339 786 341
rect 788 339 819 341
rect 821 339 822 341
rect 85 338 822 339
rect 5 333 6 335
rect 8 333 9 335
rect 5 331 9 333
rect 99 333 103 334
rect 99 331 100 333
rect 102 331 103 333
rect 99 327 103 331
rect 305 333 481 334
rect 305 331 306 333
rect 308 331 481 333
rect 305 330 478 331
rect 237 329 301 330
rect 237 327 238 329
rect 240 327 298 329
rect 300 327 301 329
rect 477 329 478 330
rect 480 329 481 331
rect 537 333 600 334
rect 537 331 538 333
rect 540 331 597 333
rect 599 331 600 333
rect 537 330 600 331
rect 637 333 641 334
rect 637 331 638 333
rect 640 331 641 333
rect 477 328 481 329
rect 605 328 609 329
rect 99 326 109 327
rect 237 326 301 327
rect 605 326 606 328
rect 608 326 609 328
rect 5 325 9 326
rect 5 323 6 325
rect 8 323 9 325
rect 99 324 106 326
rect 108 324 109 326
rect 99 323 109 324
rect 205 325 209 326
rect 205 323 206 325
rect 208 323 209 325
rect 5 297 9 323
rect 28 310 32 311
rect 28 308 29 310
rect 31 308 32 310
rect 28 304 32 308
rect 28 302 29 304
rect 31 302 32 304
rect 28 301 32 302
rect 105 305 109 323
rect 137 322 141 323
rect 137 320 138 322
rect 140 320 141 322
rect 137 315 141 320
rect 137 313 138 315
rect 140 313 141 315
rect 137 311 141 313
rect 205 313 209 323
rect 306 325 310 326
rect 306 323 307 325
rect 309 323 310 325
rect 306 322 310 323
rect 337 325 341 326
rect 337 323 338 325
rect 340 323 341 325
rect 337 320 341 323
rect 385 325 409 326
rect 385 323 386 325
rect 388 323 406 325
rect 408 323 409 325
rect 385 322 409 323
rect 437 325 441 326
rect 437 323 438 325
rect 440 323 441 325
rect 337 318 338 320
rect 340 318 341 320
rect 337 317 341 318
rect 437 321 441 323
rect 437 319 438 321
rect 440 319 441 321
rect 437 317 441 319
rect 585 325 589 326
rect 605 325 609 326
rect 637 328 641 331
rect 637 326 638 328
rect 640 326 641 328
rect 585 323 586 325
rect 588 323 589 325
rect 585 313 589 323
rect 637 319 641 326
rect 685 325 689 326
rect 685 323 686 325
rect 688 323 689 325
rect 205 309 589 313
rect 685 305 689 323
rect 705 325 709 326
rect 705 323 706 325
rect 708 323 709 325
rect 705 322 709 323
rect 785 325 789 326
rect 785 323 786 325
rect 788 323 789 325
rect 105 301 689 305
rect 728 310 732 311
rect 728 308 729 310
rect 731 308 732 310
rect 728 304 732 308
rect 728 302 729 304
rect 731 302 732 304
rect 728 301 732 302
rect 785 297 789 323
rect 5 293 789 297
rect 337 288 704 289
rect 337 286 338 288
rect 340 286 701 288
rect 703 286 704 288
rect 337 285 704 286
rect 113 277 804 281
rect 113 264 117 277
rect 113 262 114 264
rect 116 262 117 264
rect 113 261 117 262
rect 198 272 202 273
rect 198 270 199 272
rect 201 270 202 272
rect 198 263 202 270
rect 198 261 199 263
rect 201 261 202 263
rect 298 272 302 273
rect 298 270 299 272
rect 301 270 302 272
rect 298 264 302 270
rect 298 262 299 264
rect 301 262 302 264
rect 298 261 302 262
rect 313 264 317 277
rect 313 262 314 264
rect 316 262 317 264
rect 313 261 317 262
rect 495 264 504 265
rect 495 262 496 264
rect 498 262 501 264
rect 503 262 504 264
rect 495 261 504 262
rect 515 264 519 277
rect 515 262 516 264
rect 518 262 519 264
rect 515 261 519 262
rect 700 272 704 273
rect 700 270 701 272
rect 703 270 704 272
rect 700 264 704 270
rect 700 262 701 264
rect 703 262 704 264
rect 700 261 704 262
rect 715 264 719 277
rect 715 262 716 264
rect 718 262 719 264
rect 715 261 719 262
rect 198 260 202 261
rect 21 256 194 257
rect 21 254 22 256
rect 24 254 191 256
rect 193 254 194 256
rect 21 253 194 254
rect 221 256 394 257
rect 221 254 222 256
rect 224 254 391 256
rect 393 254 394 256
rect 221 253 394 254
rect 423 256 600 257
rect 423 254 424 256
rect 426 254 593 256
rect 595 254 597 256
rect 599 254 600 256
rect 423 253 600 254
rect 623 256 796 257
rect 623 254 624 256
rect 626 254 787 256
rect 789 254 793 256
rect 795 254 796 256
rect 623 253 796 254
rect 13 247 719 248
rect 13 245 14 247
rect 16 245 114 247
rect 116 245 214 247
rect 216 245 314 247
rect 316 245 416 247
rect 418 245 516 247
rect 518 245 616 247
rect 618 245 716 247
rect 718 245 719 247
rect 13 244 719 245
rect 61 239 66 240
rect 61 237 63 239
rect 65 237 66 239
rect 61 236 66 237
rect 98 239 102 240
rect 98 237 99 239
rect 101 237 102 239
rect 61 211 65 236
rect 98 235 102 237
rect 98 233 99 235
rect 101 233 102 235
rect 98 232 102 233
rect 162 239 166 240
rect 162 237 163 239
rect 165 237 166 239
rect 162 211 166 237
rect 262 239 266 240
rect 262 237 263 239
rect 265 237 266 239
rect 262 222 266 237
rect 262 220 263 222
rect 265 220 266 222
rect 262 219 266 220
rect 362 239 366 240
rect 362 237 363 239
rect 365 237 366 239
rect 61 207 102 211
rect 162 207 301 211
rect 98 205 102 207
rect 98 203 99 205
rect 101 203 102 205
rect 297 206 301 207
rect 297 204 298 206
rect 300 204 301 206
rect 362 209 366 237
rect 400 239 404 240
rect 400 237 401 239
rect 403 237 404 239
rect 400 232 404 237
rect 464 239 468 240
rect 464 237 465 239
rect 467 237 468 239
rect 464 235 468 237
rect 400 230 401 232
rect 403 230 404 232
rect 463 231 468 235
rect 400 223 404 230
rect 464 229 468 231
rect 564 239 568 240
rect 564 237 565 239
rect 567 237 568 239
rect 464 228 504 229
rect 464 226 501 228
rect 503 226 504 228
rect 464 225 504 226
rect 564 228 568 237
rect 564 226 565 228
rect 567 226 568 228
rect 564 225 568 226
rect 664 239 668 240
rect 664 237 665 239
rect 667 237 668 239
rect 664 220 668 237
rect 664 218 665 220
rect 667 218 668 220
rect 764 239 768 240
rect 764 237 765 239
rect 767 237 768 239
rect 764 221 768 237
rect 764 219 765 221
rect 767 219 768 221
rect 764 218 768 219
rect 664 217 668 218
rect 800 209 804 277
rect 362 208 396 209
rect 362 206 393 208
rect 395 206 396 208
rect 362 205 396 206
rect 400 208 804 209
rect 400 206 401 208
rect 403 206 804 208
rect 400 205 804 206
rect 297 203 301 204
rect 98 202 102 203
rect 13 197 719 198
rect 13 195 14 197
rect 16 195 114 197
rect 116 195 214 197
rect 216 195 314 197
rect 316 195 416 197
rect 418 195 516 197
rect 518 195 616 197
rect 618 195 716 197
rect 718 195 719 197
rect 13 194 719 195
rect 800 190 804 205
rect 810 221 814 222
rect 810 219 811 221
rect 813 219 814 221
rect 810 191 814 219
rect 121 189 297 190
rect 121 187 122 189
rect 124 187 294 189
rect 296 187 297 189
rect 121 186 297 187
rect 321 189 404 190
rect 321 187 322 189
rect 324 187 401 189
rect 403 187 404 189
rect 321 186 404 187
rect 495 189 504 190
rect 495 187 496 189
rect 498 187 501 189
rect 503 187 504 189
rect 495 186 504 187
rect 523 189 703 190
rect 523 187 524 189
rect 526 187 696 189
rect 698 187 700 189
rect 702 187 703 189
rect 523 186 703 187
rect 723 189 806 190
rect 723 187 724 189
rect 726 187 806 189
rect 810 189 811 191
rect 813 189 814 191
rect 810 188 814 189
rect 723 186 806 187
rect 13 181 204 182
rect 13 179 14 181
rect 16 179 194 181
rect 196 179 201 181
rect 203 179 204 181
rect 13 178 204 179
rect 213 181 396 182
rect 213 179 214 181
rect 216 179 393 181
rect 395 179 396 181
rect 213 178 396 179
rect 415 181 604 182
rect 415 179 416 181
rect 418 179 596 181
rect 598 179 601 181
rect 603 179 604 181
rect 415 178 604 179
rect 615 181 798 182
rect 615 179 616 181
rect 618 179 795 181
rect 797 179 798 181
rect 615 178 798 179
rect 61 171 65 172
rect 61 169 62 171
rect 64 169 65 171
rect 61 157 65 169
rect 170 166 201 167
rect 170 164 171 166
rect 173 164 198 166
rect 200 164 201 166
rect 170 163 201 164
rect 270 166 301 167
rect 270 164 271 166
rect 273 164 298 166
rect 300 164 301 166
rect 270 163 301 164
rect 370 166 404 167
rect 370 164 371 166
rect 373 164 401 166
rect 403 164 404 166
rect 370 163 404 164
rect 472 166 476 167
rect 472 164 473 166
rect 475 164 476 166
rect 472 157 476 164
rect 61 156 97 157
rect 61 154 94 156
rect 96 154 97 156
rect 61 153 97 154
rect 393 153 476 157
rect 572 166 576 167
rect 572 164 573 166
rect 575 164 576 166
rect 572 156 576 164
rect 672 166 704 167
rect 672 164 673 166
rect 675 164 701 166
rect 703 164 704 166
rect 672 163 704 164
rect 772 166 776 167
rect 772 164 773 166
rect 775 164 776 166
rect 572 154 573 156
rect 575 154 576 156
rect 572 153 576 154
rect 772 156 776 164
rect 772 154 773 156
rect 775 154 776 156
rect 772 153 776 154
rect 393 149 397 153
rect 13 145 397 149
rect 13 119 17 145
rect 197 140 317 141
rect 197 138 198 140
rect 200 138 317 140
rect 13 117 14 119
rect 16 117 17 119
rect 13 116 17 117
rect 93 137 97 138
rect 93 135 94 137
rect 96 135 97 137
rect 93 119 97 135
rect 93 117 94 119
rect 96 117 97 119
rect 93 116 97 117
rect 197 137 317 138
rect 197 119 201 137
rect 261 130 265 131
rect 261 128 262 130
rect 264 128 265 130
rect 261 123 265 128
rect 261 121 262 123
rect 264 121 265 123
rect 261 120 265 121
rect 197 117 198 119
rect 200 117 201 119
rect 197 116 201 117
rect 293 119 301 120
rect 293 117 294 119
rect 296 117 298 119
rect 300 117 301 119
rect 293 116 301 117
rect 313 119 317 137
rect 313 117 314 119
rect 316 117 317 119
rect 313 116 317 117
rect 393 119 397 145
rect 393 117 394 119
rect 396 117 397 119
rect 393 116 397 117
rect 415 145 798 149
rect 415 119 419 145
rect 495 140 619 141
rect 495 138 496 140
rect 498 138 619 140
rect 495 137 619 138
rect 415 117 416 119
rect 418 117 419 119
rect 415 116 419 117
rect 463 123 467 124
rect 463 121 464 123
rect 466 121 467 123
rect 61 115 65 116
rect 61 113 62 115
rect 64 113 65 115
rect 61 102 65 113
rect 121 111 297 112
rect 121 109 122 111
rect 124 109 294 111
rect 296 109 297 111
rect 121 108 297 109
rect 349 111 365 112
rect 349 109 350 111
rect 352 109 362 111
rect 364 109 365 111
rect 349 108 365 109
rect 463 111 467 121
rect 495 119 499 137
rect 495 117 496 119
rect 498 117 499 119
rect 495 116 499 117
rect 503 132 507 133
rect 503 130 504 132
rect 506 130 507 132
rect 463 109 464 111
rect 466 109 467 111
rect 463 108 467 109
rect 503 104 507 130
rect 563 132 607 133
rect 563 130 604 132
rect 606 130 607 132
rect 563 128 564 130
rect 566 129 607 130
rect 566 128 567 129
rect 563 126 567 128
rect 615 120 619 137
rect 700 138 704 139
rect 700 136 701 138
rect 703 136 704 138
rect 615 118 616 120
rect 618 118 619 120
rect 663 130 667 131
rect 663 128 664 130
rect 666 128 667 130
rect 663 122 667 128
rect 663 120 664 122
rect 666 120 667 122
rect 663 119 667 120
rect 700 119 704 136
rect 615 117 619 118
rect 700 117 701 119
rect 703 117 704 119
rect 700 116 704 117
rect 794 119 798 145
rect 794 117 795 119
rect 797 117 798 119
rect 794 116 798 117
rect 523 112 696 113
rect 523 110 524 112
rect 526 110 693 112
rect 695 110 696 112
rect 523 109 696 110
rect 802 107 806 186
rect 810 156 814 157
rect 810 154 811 156
rect 813 154 814 156
rect 810 119 814 154
rect 810 117 811 119
rect 813 117 814 119
rect 810 116 814 117
rect 723 106 806 107
rect 723 104 724 106
rect 726 104 806 106
rect 61 100 62 102
rect 64 100 65 102
rect 161 103 209 104
rect 161 101 162 103
rect 164 101 206 103
rect 208 101 209 103
rect 161 100 209 101
rect 221 103 603 104
rect 723 103 806 104
rect 221 101 222 103
rect 224 101 600 103
rect 602 101 603 103
rect 221 100 603 101
rect 61 99 65 100
rect 763 98 767 99
rect 763 96 764 98
rect 766 96 767 98
rect 22 94 728 95
rect 22 92 23 94
rect 25 92 122 94
rect 124 92 222 94
rect 224 92 322 94
rect 324 92 424 94
rect 426 92 525 94
rect 527 92 625 94
rect 627 92 725 94
rect 727 92 728 94
rect 22 91 728 92
rect 5 88 9 89
rect 5 86 6 88
rect 8 86 9 88
rect 5 37 9 86
rect 401 86 607 87
rect 401 84 402 86
rect 404 84 604 86
rect 606 84 607 86
rect 401 83 607 84
rect 763 78 767 96
rect 77 74 767 78
rect 77 54 81 74
rect 177 69 604 70
rect 177 67 464 69
rect 466 67 604 69
rect 177 66 604 67
rect 177 62 181 66
rect 600 62 604 66
rect 177 60 178 62
rect 180 60 181 62
rect 177 59 181 60
rect 277 61 504 62
rect 277 59 278 61
rect 280 59 501 61
rect 503 59 504 61
rect 600 60 601 62
rect 603 60 604 62
rect 600 59 604 60
rect 701 61 705 74
rect 701 59 702 61
rect 704 59 705 61
rect 277 58 504 59
rect 701 58 705 59
rect 77 52 78 54
rect 80 52 81 54
rect 77 51 81 52
rect 85 53 822 54
rect 85 51 86 53
rect 88 51 186 53
rect 188 51 286 53
rect 288 51 386 53
rect 388 51 486 53
rect 488 51 586 53
rect 588 51 686 53
rect 688 51 786 53
rect 788 51 819 53
rect 821 51 822 53
rect 85 50 822 51
rect 205 45 209 46
rect 137 44 141 45
rect 137 42 138 44
rect 140 42 141 44
rect 137 41 141 42
rect 205 43 206 45
rect 208 43 209 45
rect 5 35 6 37
rect 8 35 9 37
rect 5 9 9 35
rect 105 38 109 39
rect 105 36 106 38
rect 108 36 109 38
rect 28 22 32 23
rect 28 20 29 22
rect 31 20 32 22
rect 28 19 32 20
rect 105 17 109 36
rect 205 37 209 43
rect 301 45 481 46
rect 301 43 302 45
rect 304 43 306 45
rect 308 43 481 45
rect 301 42 478 43
rect 237 41 241 42
rect 237 39 238 41
rect 240 39 241 41
rect 477 41 478 42
rect 480 41 481 43
rect 505 45 609 46
rect 505 43 506 45
rect 508 43 609 45
rect 505 42 609 43
rect 477 40 481 41
rect 237 38 241 39
rect 605 38 609 42
rect 205 35 206 37
rect 208 35 209 37
rect 385 37 409 38
rect 385 35 386 37
rect 388 35 402 37
rect 404 35 406 37
rect 408 35 409 37
rect 585 37 589 38
rect 585 35 586 37
rect 588 35 589 37
rect 205 25 209 35
rect 337 34 341 35
rect 385 34 409 35
rect 337 32 338 34
rect 340 32 341 34
rect 337 30 341 32
rect 437 33 441 35
rect 437 31 438 33
rect 440 31 441 33
rect 437 30 441 31
rect 537 33 541 35
rect 537 31 538 33
rect 540 31 541 33
rect 537 30 541 31
rect 585 25 589 35
rect 605 37 667 38
rect 605 35 664 37
rect 666 35 667 37
rect 605 34 667 35
rect 685 37 689 38
rect 685 35 686 37
rect 688 35 689 37
rect 785 37 789 38
rect 785 35 786 37
rect 788 35 789 37
rect 205 21 589 25
rect 637 27 641 28
rect 637 25 638 27
rect 640 25 641 27
rect 637 23 641 25
rect 685 17 689 35
rect 737 33 741 35
rect 737 31 738 33
rect 740 31 741 33
rect 737 30 741 31
rect 105 16 689 17
rect 105 14 350 16
rect 352 14 689 16
rect 105 13 689 14
rect 785 9 789 35
rect 5 5 789 9
rect 94 -3 98 -2
rect 94 -5 95 -3
rect 97 -5 98 -3
rect 67 -54 72 -52
rect 67 -56 68 -54
rect 70 -56 72 -54
rect 67 -58 72 -56
rect 94 -53 98 -5
rect 94 -55 95 -53
rect 97 -55 98 -53
rect 94 -57 98 -55
rect 172 -54 178 -52
rect 172 -56 174 -54
rect 176 -56 178 -54
rect 172 -58 178 -56
rect 200 -54 204 -52
rect 200 -56 201 -54
rect 203 -56 204 -54
rect 200 -57 204 -56
rect 279 -54 284 -52
rect 279 -56 280 -54
rect 282 -56 284 -54
rect 306 -53 310 -52
rect 306 -55 307 -53
rect 309 -55 310 -53
rect 306 -56 310 -55
rect 385 -54 390 -52
rect 385 -56 386 -54
rect 388 -56 390 -54
rect 279 -58 284 -56
rect 385 -58 390 -56
rect 412 -54 416 -52
rect 412 -56 413 -54
rect 415 -56 416 -54
rect 412 -57 416 -56
rect 489 -55 496 -52
rect 489 -57 491 -55
rect 493 -57 496 -55
rect 489 -58 496 -57
rect 518 -54 522 -52
rect 518 -56 519 -54
rect 521 -56 522 -54
rect 518 -58 522 -56
rect 596 -54 602 -52
rect 596 -56 598 -54
rect 600 -56 602 -54
rect 596 -58 602 -56
rect 624 -54 628 -52
rect 624 -56 625 -54
rect 627 -56 628 -54
rect 624 -58 628 -56
rect 700 -54 708 -52
rect 700 -56 702 -54
rect 704 -56 708 -54
rect 700 -58 708 -56
rect 730 -55 734 -52
rect 730 -57 731 -55
rect 733 -57 734 -55
rect 730 -58 734 -57
rect 807 -54 814 -52
rect 807 -56 809 -54
rect 811 -56 814 -54
rect 807 -58 814 -56
rect 914 -54 920 -52
rect 914 -56 916 -54
rect 918 -56 920 -54
rect 914 -58 920 -56
rect -12 -62 -7 -61
rect -12 -64 -11 -62
rect -9 -64 -7 -62
rect -12 -66 -7 -64
rect 59 -78 912 -77
rect 59 -80 61 -78
rect 63 -80 167 -78
rect 169 -80 273 -78
rect 275 -80 379 -78
rect 381 -80 485 -78
rect 487 -80 591 -78
rect 593 -80 697 -78
rect 699 -80 803 -78
rect 805 -80 909 -78
rect 911 -80 912 -78
rect 59 -81 912 -80
<< alu3 >>
rect 308 1166 318 1167
rect 284 1163 288 1165
rect 284 1161 285 1163
rect 287 1161 288 1163
rect 209 1159 213 1160
rect 284 1159 288 1161
rect 308 1164 315 1166
rect 317 1164 318 1166
rect 308 1163 318 1164
rect 347 1163 373 1164
rect 209 1157 210 1159
rect 212 1157 213 1159
rect 209 1112 213 1157
rect 209 1108 242 1112
rect 144 1107 205 1108
rect 144 1105 145 1107
rect 147 1105 202 1107
rect 204 1105 205 1107
rect 144 1104 205 1105
rect 72 1085 167 1086
rect 72 1083 164 1085
rect 166 1083 167 1085
rect 72 1082 167 1083
rect 50 1013 54 1015
rect 50 1011 51 1013
rect 53 1011 54 1013
rect 50 985 54 1011
rect 50 983 51 985
rect 53 983 54 985
rect 50 982 54 983
rect 72 829 76 1082
rect 173 1071 233 1072
rect 173 1069 174 1071
rect 176 1069 230 1071
rect 232 1069 233 1071
rect 173 1068 233 1069
rect 238 1056 242 1108
rect 80 1055 242 1056
rect 80 1053 81 1055
rect 83 1053 242 1055
rect 80 1052 242 1053
rect 80 928 84 929
rect 80 926 81 928
rect 83 926 84 928
rect 80 925 84 926
rect 80 924 108 925
rect 80 922 105 924
rect 107 922 108 924
rect 80 921 108 922
rect 112 839 116 1052
rect 156 1037 160 1038
rect 156 1035 157 1037
rect 159 1035 160 1037
rect 133 1028 137 1029
rect 133 1026 134 1028
rect 136 1026 137 1028
rect 120 924 124 925
rect 120 922 121 924
rect 123 922 124 924
rect 120 901 124 922
rect 120 899 121 901
rect 123 899 124 901
rect 120 898 124 899
rect 112 837 113 839
rect 115 837 116 839
rect 112 836 116 837
rect 133 829 137 1026
rect 72 825 137 829
rect 148 963 152 964
rect 148 961 149 963
rect 151 961 152 963
rect 148 949 152 961
rect 148 947 149 949
rect 151 947 152 949
rect 148 891 152 947
rect 148 889 149 891
rect 151 889 152 891
rect 72 778 76 825
rect 148 820 152 889
rect 156 883 160 1035
rect 156 881 157 883
rect 159 881 160 883
rect 156 880 160 881
rect 180 883 184 1052
rect 308 1048 312 1163
rect 347 1161 348 1163
rect 350 1161 373 1163
rect 347 1160 373 1161
rect 212 1047 216 1048
rect 212 1045 213 1047
rect 215 1045 216 1047
rect 200 934 204 937
rect 200 932 201 934
rect 203 932 204 934
rect 200 931 204 932
rect 212 925 216 1045
rect 220 1047 312 1048
rect 220 1045 221 1047
rect 223 1045 312 1047
rect 220 1044 312 1045
rect 271 993 275 994
rect 271 991 272 993
rect 274 991 275 993
rect 271 951 275 991
rect 308 951 312 1044
rect 271 950 312 951
rect 271 948 272 950
rect 274 948 309 950
rect 311 948 312 950
rect 271 947 312 948
rect 336 1107 340 1108
rect 336 1105 337 1107
rect 339 1105 340 1107
rect 336 1054 340 1105
rect 336 1052 337 1054
rect 339 1052 340 1054
rect 212 924 273 925
rect 212 922 270 924
rect 272 922 273 924
rect 212 921 273 922
rect 180 881 181 883
rect 183 881 184 883
rect 180 839 184 881
rect 220 875 258 876
rect 220 873 221 875
rect 223 873 255 875
rect 257 873 258 875
rect 220 872 258 873
rect 203 852 210 853
rect 203 850 204 852
rect 206 850 210 852
rect 203 849 210 850
rect 180 837 181 839
rect 183 837 184 839
rect 180 836 184 837
rect 206 820 210 849
rect 269 839 273 921
rect 336 892 340 1052
rect 344 1062 348 1063
rect 344 1060 345 1062
rect 347 1060 348 1062
rect 344 901 348 1060
rect 369 1013 373 1160
rect 660 1162 664 1164
rect 660 1160 661 1162
rect 663 1160 664 1162
rect 660 1158 664 1160
rect 555 1107 743 1108
rect 555 1105 556 1107
rect 558 1105 740 1107
rect 742 1105 743 1107
rect 555 1104 743 1105
rect 764 1093 826 1094
rect 764 1091 766 1093
rect 768 1091 826 1093
rect 764 1090 826 1091
rect 573 1081 577 1082
rect 573 1079 574 1081
rect 576 1079 577 1081
rect 369 1011 370 1013
rect 372 1011 373 1013
rect 369 1010 373 1011
rect 407 1052 433 1053
rect 407 1051 567 1052
rect 407 1049 564 1051
rect 566 1049 567 1051
rect 407 1048 567 1049
rect 344 899 345 901
rect 347 899 348 901
rect 344 898 348 899
rect 324 891 340 892
rect 324 889 325 891
rect 327 889 340 891
rect 324 888 340 889
rect 269 837 270 839
rect 272 837 273 839
rect 269 836 273 837
rect 116 819 201 820
rect 116 817 198 819
rect 200 817 201 819
rect 116 816 201 817
rect 206 819 284 820
rect 206 817 281 819
rect 283 817 284 819
rect 206 816 284 817
rect 116 797 120 816
rect 116 795 117 797
rect 119 795 120 797
rect 116 794 120 795
rect 275 798 279 799
rect 275 796 276 798
rect 278 796 279 798
rect 72 777 100 778
rect 72 775 97 777
rect 99 775 100 777
rect 72 774 100 775
rect 124 747 266 748
rect 124 745 125 747
rect 127 745 263 747
rect 265 745 266 747
rect 124 744 266 745
rect 50 722 54 724
rect 31 719 35 721
rect 31 717 32 719
rect 34 717 35 719
rect 31 692 35 717
rect 50 720 51 722
rect 53 720 54 722
rect 50 703 54 720
rect 50 701 51 703
rect 53 701 54 703
rect 50 700 54 701
rect 31 690 32 692
rect 34 690 35 692
rect 31 689 35 690
rect 275 683 279 796
rect 308 731 312 733
rect 308 729 309 731
rect 311 729 312 731
rect 308 727 312 729
rect 275 681 276 683
rect 278 681 279 683
rect 275 680 279 681
rect 184 632 373 633
rect 184 630 370 632
rect 372 630 373 632
rect 184 629 373 630
rect 184 623 188 629
rect 184 621 185 623
rect 187 621 188 623
rect 184 598 188 621
rect 184 596 185 598
rect 187 596 188 598
rect 31 589 35 596
rect 184 595 188 596
rect 246 623 381 624
rect 246 621 247 623
rect 249 621 378 623
rect 380 621 381 623
rect 246 620 381 621
rect 31 587 32 589
rect 34 587 35 589
rect 20 582 24 584
rect 20 580 21 582
rect 23 580 24 582
rect 20 554 24 580
rect 20 552 21 554
rect 23 552 24 554
rect 20 549 24 552
rect 31 552 35 587
rect 31 550 32 552
rect 34 550 35 552
rect 31 548 35 550
rect 50 581 54 583
rect 50 579 51 581
rect 53 579 54 581
rect 50 553 54 579
rect 246 577 250 620
rect 407 608 411 1048
rect 573 1036 577 1079
rect 442 1035 577 1036
rect 442 1033 443 1035
rect 445 1033 574 1035
rect 576 1033 577 1035
rect 442 1032 577 1033
rect 635 1060 639 1061
rect 635 1058 636 1060
rect 638 1058 639 1060
rect 635 1035 639 1058
rect 635 1033 636 1035
rect 638 1033 639 1035
rect 635 1027 639 1033
rect 450 1026 639 1027
rect 450 1024 451 1026
rect 453 1024 639 1026
rect 450 1023 639 1024
rect 544 975 548 976
rect 544 973 545 975
rect 547 973 548 975
rect 511 926 515 929
rect 511 924 512 926
rect 514 924 515 926
rect 511 922 515 924
rect 544 860 548 973
rect 723 881 751 882
rect 723 879 724 881
rect 726 879 751 881
rect 723 878 751 879
rect 695 867 699 869
rect 695 865 696 867
rect 698 865 699 867
rect 695 862 699 865
rect 544 858 545 860
rect 547 858 548 860
rect 544 857 548 858
rect 703 861 707 862
rect 703 859 704 861
rect 706 859 707 861
rect 703 840 707 859
rect 539 839 617 840
rect 539 837 540 839
rect 542 837 617 839
rect 539 836 617 837
rect 622 839 707 840
rect 622 837 623 839
rect 625 837 707 839
rect 622 836 707 837
rect 550 819 554 820
rect 550 817 551 819
rect 553 817 554 819
rect 483 767 499 768
rect 483 765 496 767
rect 498 765 499 767
rect 483 764 499 765
rect 475 757 479 758
rect 475 755 476 757
rect 478 755 479 757
rect 256 607 411 608
rect 256 605 257 607
rect 259 605 411 607
rect 256 604 411 605
rect 450 645 454 646
rect 450 643 451 645
rect 453 643 454 645
rect 246 575 247 577
rect 249 575 250 577
rect 246 574 250 575
rect 50 551 51 553
rect 53 551 54 553
rect 50 549 54 551
rect 80 551 268 552
rect 80 549 81 551
rect 83 549 265 551
rect 267 549 268 551
rect 80 548 268 549
rect 159 497 163 500
rect 159 495 160 497
rect 162 495 163 497
rect 159 493 163 495
rect 450 496 454 643
rect 475 596 479 755
rect 475 594 476 596
rect 478 594 479 596
rect 475 593 479 594
rect 483 604 487 764
rect 550 735 554 817
rect 613 807 617 836
rect 639 819 643 820
rect 639 817 640 819
rect 642 817 643 819
rect 613 806 620 807
rect 613 804 617 806
rect 619 804 620 806
rect 613 803 620 804
rect 565 783 603 784
rect 565 781 566 783
rect 568 781 600 783
rect 602 781 603 783
rect 565 780 603 781
rect 639 775 643 817
rect 639 773 640 775
rect 642 773 643 775
rect 550 734 611 735
rect 550 732 551 734
rect 553 732 611 734
rect 550 731 611 732
rect 483 602 484 604
rect 486 602 487 604
rect 483 551 487 602
rect 483 549 484 551
rect 486 549 487 551
rect 483 548 487 549
rect 511 708 552 709
rect 511 706 512 708
rect 514 706 549 708
rect 551 706 552 708
rect 511 705 552 706
rect 511 612 515 705
rect 548 665 552 705
rect 548 663 549 665
rect 551 663 552 665
rect 548 662 552 663
rect 511 611 603 612
rect 511 609 600 611
rect 602 609 603 611
rect 511 608 603 609
rect 607 611 611 731
rect 619 723 623 726
rect 619 721 620 723
rect 622 721 623 723
rect 619 719 623 721
rect 607 609 608 611
rect 610 609 611 611
rect 607 608 611 609
rect 450 495 476 496
rect 450 493 473 495
rect 475 493 476 495
rect 511 493 515 608
rect 639 604 643 773
rect 663 775 667 776
rect 663 773 664 775
rect 666 773 667 775
rect 663 621 667 773
rect 671 767 675 836
rect 747 831 751 878
rect 671 765 672 767
rect 674 765 675 767
rect 671 709 675 765
rect 671 707 672 709
rect 674 707 675 709
rect 671 695 675 707
rect 671 693 672 695
rect 674 693 675 695
rect 671 692 675 693
rect 686 827 751 831
rect 686 630 690 827
rect 707 819 711 820
rect 707 817 708 819
rect 710 817 711 819
rect 699 757 703 758
rect 699 755 700 757
rect 702 755 703 757
rect 699 734 703 755
rect 699 732 700 734
rect 702 732 703 734
rect 699 731 703 732
rect 686 628 687 630
rect 689 628 690 630
rect 686 627 690 628
rect 663 619 664 621
rect 666 619 667 621
rect 663 618 667 619
rect 707 604 711 817
rect 715 734 743 735
rect 715 732 716 734
rect 718 732 743 734
rect 715 731 743 732
rect 739 730 743 731
rect 739 728 740 730
rect 742 728 743 730
rect 739 727 743 728
rect 581 603 743 604
rect 581 601 740 603
rect 742 601 743 603
rect 581 600 743 601
rect 581 548 585 600
rect 590 587 650 588
rect 590 585 591 587
rect 593 585 647 587
rect 649 585 650 587
rect 590 584 650 585
rect 747 574 751 827
rect 656 573 751 574
rect 656 571 657 573
rect 659 571 751 573
rect 656 570 751 571
rect 618 551 679 552
rect 618 549 619 551
rect 621 549 676 551
rect 678 549 679 551
rect 618 548 679 549
rect 581 544 614 548
rect 610 499 614 544
rect 610 497 611 499
rect 613 497 614 499
rect 450 492 476 493
rect 505 492 515 493
rect 505 490 506 492
rect 508 490 515 492
rect 535 495 539 497
rect 610 496 614 497
rect 535 493 536 495
rect 538 493 539 495
rect 535 491 539 493
rect 505 489 515 490
rect 705 457 709 458
rect 705 455 706 457
rect 708 455 709 457
rect 705 454 709 455
rect 822 448 826 1090
rect 689 447 826 448
rect 689 445 691 447
rect 693 445 826 447
rect 689 444 826 445
rect 605 435 635 436
rect 605 433 630 435
rect 632 433 635 435
rect 605 432 635 433
rect 500 422 504 423
rect 500 420 501 422
rect 503 420 504 422
rect 266 382 271 383
rect 266 380 267 382
rect 269 380 271 382
rect 266 379 271 380
rect 99 378 103 379
rect 99 376 100 378
rect 102 376 103 378
rect 99 333 103 376
rect 201 374 205 375
rect 201 372 202 374
rect 204 372 205 374
rect 201 349 205 372
rect 201 347 202 349
rect 204 347 205 349
rect 201 346 205 347
rect 500 349 504 420
rect 500 347 501 349
rect 503 347 504 349
rect 500 346 504 347
rect 99 331 100 333
rect 102 331 103 333
rect 99 330 103 331
rect 198 334 441 338
rect 137 315 141 316
rect 137 313 138 315
rect 140 313 141 315
rect 28 304 32 305
rect 28 302 29 304
rect 31 302 32 304
rect 28 285 32 302
rect 28 281 102 285
rect 98 235 102 281
rect 137 252 141 313
rect 198 272 202 334
rect 297 329 302 330
rect 297 327 298 329
rect 300 327 302 329
rect 297 326 302 327
rect 198 270 199 272
rect 201 270 202 272
rect 198 269 202 270
rect 298 272 302 326
rect 306 325 310 326
rect 306 323 307 325
rect 309 323 310 325
rect 306 322 310 323
rect 405 325 409 326
rect 405 323 406 325
rect 408 323 409 325
rect 405 322 409 323
rect 437 325 441 334
rect 437 323 438 325
rect 440 323 441 325
rect 437 322 441 323
rect 596 333 600 334
rect 596 331 597 333
rect 599 331 600 333
rect 337 320 341 321
rect 337 318 338 320
rect 340 318 341 320
rect 337 288 341 318
rect 337 286 338 288
rect 340 286 341 288
rect 337 285 341 286
rect 298 270 299 272
rect 301 270 302 272
rect 298 269 302 270
rect 495 264 499 265
rect 495 262 496 264
rect 498 262 499 264
rect 495 252 499 262
rect 596 256 600 331
rect 605 328 609 432
rect 818 341 822 342
rect 818 339 819 341
rect 821 339 822 341
rect 605 326 606 328
rect 608 326 609 328
rect 605 325 609 326
rect 637 328 641 329
rect 637 326 638 328
rect 640 326 641 328
rect 596 254 597 256
rect 599 254 600 256
rect 596 253 600 254
rect 137 248 499 252
rect 637 237 641 326
rect 705 325 709 326
rect 705 323 706 325
rect 708 323 709 325
rect 705 322 709 323
rect 728 304 790 305
rect 728 302 729 304
rect 731 302 790 304
rect 728 301 790 302
rect 700 288 704 289
rect 700 286 701 288
rect 703 286 704 288
rect 700 272 704 286
rect 700 270 701 272
rect 703 270 704 272
rect 700 269 704 270
rect 786 256 790 301
rect 786 254 787 256
rect 789 254 790 256
rect 786 253 790 254
rect 98 233 99 235
rect 101 233 102 235
rect 478 233 641 237
rect 98 232 102 233
rect 400 232 404 233
rect 400 230 401 232
rect 403 230 404 232
rect 400 227 404 230
rect 478 227 482 233
rect 400 223 482 227
rect 500 228 504 229
rect 500 226 501 228
rect 503 226 504 228
rect 200 222 266 223
rect 200 220 263 222
rect 265 220 266 222
rect 200 219 266 220
rect 200 181 204 219
rect 400 208 404 209
rect 400 206 401 208
rect 403 206 404 208
rect 400 189 404 206
rect 400 187 401 189
rect 403 187 404 189
rect 400 186 404 187
rect 500 189 504 226
rect 564 228 703 229
rect 564 226 565 228
rect 567 226 703 228
rect 564 225 703 226
rect 500 187 501 189
rect 503 187 504 189
rect 500 186 504 187
rect 600 220 668 221
rect 600 218 665 220
rect 667 218 668 220
rect 600 217 668 218
rect 200 179 201 181
rect 203 179 204 181
rect 200 178 204 179
rect 600 181 604 217
rect 699 189 703 225
rect 764 221 814 222
rect 764 219 765 221
rect 767 219 811 221
rect 813 219 814 221
rect 764 218 814 219
rect 699 187 700 189
rect 702 187 703 189
rect 699 186 703 187
rect 600 179 601 181
rect 603 179 604 181
rect 600 178 604 179
rect 197 166 201 167
rect 197 164 198 166
rect 200 164 201 166
rect 93 156 97 157
rect 93 154 94 156
rect 96 154 97 156
rect 93 137 97 154
rect 197 140 201 164
rect 197 138 198 140
rect 200 138 201 140
rect 197 137 201 138
rect 297 166 301 167
rect 297 164 298 166
rect 300 164 301 166
rect 93 135 94 137
rect 96 135 97 137
rect 93 134 97 135
rect 297 133 301 164
rect 400 166 499 167
rect 400 164 401 166
rect 403 164 499 166
rect 400 163 499 164
rect 495 140 499 163
rect 700 166 704 167
rect 700 164 701 166
rect 703 164 704 166
rect 495 138 496 140
rect 498 138 499 140
rect 495 137 499 138
rect 572 156 576 157
rect 572 154 573 156
rect 575 154 576 156
rect 297 132 507 133
rect 297 130 504 132
rect 506 130 507 132
rect 297 129 507 130
rect 261 123 265 124
rect 261 121 262 123
rect 264 121 265 123
rect 261 112 265 121
rect 572 120 576 154
rect 700 138 704 164
rect 772 156 814 157
rect 772 154 773 156
rect 775 154 811 156
rect 813 154 814 156
rect 772 153 814 154
rect 700 136 701 138
rect 703 136 704 138
rect 700 135 704 136
rect 293 119 576 120
rect 293 117 298 119
rect 300 117 576 119
rect 293 116 576 117
rect 603 132 607 133
rect 603 130 604 132
rect 606 130 607 132
rect 261 108 305 112
rect 205 103 209 104
rect 61 102 65 103
rect 61 100 62 102
rect 64 100 65 102
rect 61 89 65 100
rect 5 88 65 89
rect 5 86 6 88
rect 8 86 65 88
rect 5 85 65 86
rect 205 101 206 103
rect 208 101 209 103
rect 205 45 209 101
rect 137 44 141 45
rect 137 42 138 44
rect 140 42 141 44
rect 205 43 206 45
rect 208 43 209 45
rect 205 42 209 43
rect 301 45 305 108
rect 301 43 302 45
rect 304 43 305 45
rect 301 42 305 43
rect 349 111 353 112
rect 349 109 350 111
rect 352 109 353 111
rect 28 22 32 23
rect 28 20 29 22
rect 31 20 32 22
rect 28 -6 32 20
rect 137 -2 141 42
rect 94 -3 141 -2
rect 94 -5 95 -3
rect 97 -5 141 -3
rect 94 -6 141 -5
rect 237 41 241 42
rect 237 39 238 41
rect 240 39 241 41
rect -12 -10 32 -6
rect 237 -8 241 39
rect 337 34 341 35
rect 337 32 338 34
rect 340 32 341 34
rect 337 -2 341 32
rect 349 16 353 109
rect 463 111 467 112
rect 463 109 464 111
rect 466 109 467 111
rect 401 86 405 87
rect 401 84 402 86
rect 404 84 405 86
rect 401 37 405 84
rect 463 69 467 109
rect 603 86 607 130
rect 603 84 604 86
rect 606 84 607 86
rect 603 83 607 84
rect 663 122 667 124
rect 663 120 664 122
rect 666 120 667 122
rect 463 67 464 69
rect 466 67 467 69
rect 463 66 467 67
rect 401 35 402 37
rect 404 35 405 37
rect 663 37 667 120
rect 818 53 822 339
rect 818 51 819 53
rect 821 51 822 53
rect 818 50 822 51
rect 663 35 664 37
rect 666 35 667 37
rect 401 34 405 35
rect 349 14 350 16
rect 352 14 353 16
rect 349 13 353 14
rect 437 33 441 35
rect 437 31 438 33
rect 440 31 441 33
rect -12 -62 -8 -10
rect 200 -12 241 -8
rect 306 -6 341 -2
rect -12 -64 -11 -62
rect -9 -64 -8 -62
rect -12 -66 -8 -64
rect 67 -54 72 -52
rect 67 -56 68 -54
rect 70 -56 72 -54
rect 67 -112 72 -56
rect 67 -114 68 -112
rect 70 -114 72 -112
rect 67 -116 72 -114
rect 172 -54 178 -52
rect 172 -56 174 -54
rect 176 -56 178 -54
rect 172 -167 178 -56
rect 200 -54 204 -12
rect 200 -56 201 -54
rect 203 -56 204 -54
rect 200 -57 204 -56
rect 279 -54 284 -52
rect 279 -56 280 -54
rect 282 -56 284 -54
rect 306 -53 310 -6
rect 437 -8 441 31
rect 537 33 541 35
rect 663 34 667 35
rect 537 31 538 33
rect 540 31 541 33
rect 537 -7 541 31
rect 737 33 741 35
rect 737 31 738 33
rect 740 31 741 33
rect 412 -12 441 -8
rect 518 -11 541 -7
rect 637 27 641 28
rect 637 25 638 27
rect 640 25 641 27
rect 637 -8 641 25
rect 306 -55 307 -53
rect 309 -55 310 -53
rect 306 -56 310 -55
rect 385 -54 390 -52
rect 385 -56 386 -54
rect 388 -56 390 -54
rect 172 -169 174 -167
rect 176 -169 178 -167
rect 172 -171 178 -169
rect 279 -184 284 -56
rect 279 -186 281 -184
rect 283 -186 284 -184
rect 279 -187 284 -186
rect 385 -208 390 -56
rect 412 -54 416 -12
rect 412 -56 413 -54
rect 415 -56 416 -54
rect 412 -57 416 -56
rect 489 -55 496 -52
rect 489 -57 491 -55
rect 493 -57 496 -55
rect 385 -210 387 -208
rect 389 -210 390 -208
rect 385 -211 390 -210
rect 489 -278 496 -57
rect 518 -54 522 -11
rect 624 -12 641 -8
rect 737 -10 741 31
rect 518 -56 519 -54
rect 521 -56 522 -54
rect 518 -58 522 -56
rect 596 -54 602 -52
rect 596 -56 598 -54
rect 600 -56 602 -54
rect 596 -268 602 -56
rect 624 -54 628 -12
rect 730 -14 741 -10
rect 624 -56 625 -54
rect 627 -56 628 -54
rect 624 -58 628 -56
rect 700 -54 708 -52
rect 700 -56 702 -54
rect 704 -56 708 -54
rect 700 -58 708 -56
rect 730 -55 734 -14
rect 730 -57 731 -55
rect 733 -57 734 -55
rect 730 -58 734 -57
rect 807 -54 814 -52
rect 807 -56 809 -54
rect 811 -56 814 -54
rect 807 -58 814 -56
rect 914 -54 920 -52
rect 914 -56 916 -54
rect 918 -56 920 -54
rect 700 -215 706 -58
rect 807 -186 811 -58
rect 807 -188 808 -186
rect 810 -188 811 -186
rect 807 -189 811 -188
rect 700 -217 702 -215
rect 704 -217 706 -215
rect 700 -218 706 -217
rect 914 -259 920 -56
rect 914 -261 916 -259
rect 918 -261 920 -259
rect 914 -262 920 -261
rect 596 -270 598 -268
rect 600 -270 602 -268
rect 596 -271 602 -270
rect 489 -280 491 -278
rect 493 -280 496 -278
rect 489 -281 496 -280
<< alu4 >>
rect 284 1163 288 1165
rect -79 1161 285 1163
rect 287 1161 288 1163
rect -79 1159 288 1161
rect 660 1163 664 1164
rect 660 1162 1070 1163
rect 660 1160 661 1162
rect 663 1160 1070 1162
rect 660 1159 1070 1160
rect -79 -207 -75 1159
rect 660 1158 664 1159
rect -57 934 204 935
rect -57 932 201 934
rect 203 932 204 934
rect -57 931 204 932
rect -57 -183 -53 931
rect 511 926 515 927
rect 511 924 512 926
rect 514 924 1058 926
rect 511 922 1058 924
rect 695 868 699 869
rect 695 867 1033 868
rect 695 865 696 867
rect 698 865 1033 867
rect 695 864 1033 865
rect 695 862 699 864
rect 308 732 312 733
rect -42 731 312 732
rect -42 729 309 731
rect 311 729 312 731
rect -42 727 312 729
rect -42 -166 -37 727
rect 619 723 1020 724
rect 619 721 620 723
rect 622 721 1020 723
rect 619 720 1020 721
rect 619 719 623 720
rect 159 498 163 500
rect -27 497 163 498
rect -27 495 160 497
rect 162 495 163 497
rect -27 493 163 495
rect 535 495 539 496
rect 535 493 536 495
rect 538 493 991 495
rect -27 -111 -22 493
rect 535 491 991 493
rect 705 457 709 458
rect 705 455 706 457
rect 708 455 709 457
rect 405 447 695 448
rect 405 445 691 447
rect 693 445 695 447
rect 405 444 695 445
rect 266 382 310 383
rect 266 380 267 382
rect 269 380 310 382
rect 266 379 310 380
rect 306 325 310 379
rect 306 323 307 325
rect 309 323 310 325
rect 306 322 310 323
rect 405 325 409 444
rect 405 323 406 325
rect 408 323 409 325
rect 405 322 409 323
rect 705 325 709 455
rect 705 323 706 325
rect 708 323 709 325
rect 705 322 709 323
rect -27 -112 72 -111
rect -27 -114 68 -112
rect 70 -114 72 -112
rect -27 -116 72 -114
rect -42 -167 178 -166
rect -42 -169 174 -167
rect 176 -169 178 -167
rect -42 -171 178 -169
rect -57 -184 284 -183
rect -57 -186 281 -184
rect 283 -186 284 -184
rect 987 -185 991 491
rect -57 -187 284 -186
rect 807 -186 991 -185
rect 807 -188 808 -186
rect 810 -188 991 -186
rect 807 -189 991 -188
rect -79 -208 390 -207
rect -79 -210 387 -208
rect 389 -210 390 -208
rect -79 -211 390 -210
rect 1016 -214 1020 720
rect 700 -215 1020 -214
rect 700 -217 702 -215
rect 704 -217 1020 -215
rect 700 -218 1020 -217
rect 1029 -258 1033 864
rect 914 -259 1033 -258
rect 914 -261 916 -259
rect 918 -261 1033 -259
rect 914 -262 1033 -261
rect 1054 -267 1058 922
rect 596 -268 1058 -267
rect 596 -270 598 -268
rect 600 -270 1058 -268
rect 596 -271 1058 -270
rect 1066 -277 1070 1159
rect 489 -278 1070 -277
rect 489 -280 491 -278
rect 493 -280 1070 -278
rect 489 -281 1070 -280
<< ptie >>
rect 81 1183 87 1185
rect 81 1181 83 1183
rect 85 1181 87 1183
rect 81 1179 87 1181
rect 169 1183 175 1185
rect 169 1181 171 1183
rect 173 1181 175 1183
rect 169 1179 175 1181
rect 185 1183 191 1185
rect 185 1181 187 1183
rect 189 1181 191 1183
rect 185 1179 191 1181
rect 229 1183 235 1185
rect 229 1181 231 1183
rect 233 1181 235 1183
rect 229 1179 235 1181
rect 359 1183 377 1185
rect 359 1181 361 1183
rect 363 1181 373 1183
rect 375 1181 377 1183
rect 359 1179 377 1181
rect 567 1183 593 1185
rect 567 1181 569 1183
rect 571 1181 589 1183
rect 591 1181 593 1183
rect 567 1179 593 1181
rect 605 1183 611 1185
rect 605 1181 607 1183
rect 609 1181 611 1183
rect 605 1179 611 1181
rect 676 1183 694 1185
rect 676 1181 678 1183
rect 680 1181 690 1183
rect 692 1181 694 1183
rect 676 1179 694 1181
rect 700 1183 706 1185
rect 700 1181 702 1183
rect 704 1181 706 1183
rect 700 1170 706 1181
rect 117 1051 135 1053
rect 117 1049 119 1051
rect 121 1049 131 1051
rect 133 1049 135 1051
rect 117 1047 135 1049
rect 145 1051 151 1053
rect 145 1049 147 1051
rect 149 1049 151 1051
rect 145 1047 151 1049
rect 189 1051 195 1053
rect 189 1049 191 1051
rect 193 1049 195 1051
rect 189 1047 195 1049
rect 321 1051 327 1068
rect 321 1049 323 1051
rect 325 1049 327 1051
rect 321 1047 327 1049
rect 570 1051 588 1053
rect 570 1049 572 1051
rect 574 1049 584 1051
rect 586 1049 588 1051
rect 570 1047 588 1049
rect 602 1051 608 1053
rect 602 1049 604 1051
rect 606 1049 608 1051
rect 602 1047 608 1049
rect 736 1051 742 1053
rect 736 1049 738 1051
rect 740 1049 742 1051
rect 736 1047 742 1049
rect 81 1039 87 1041
rect 81 1037 83 1039
rect 85 1037 87 1039
rect 81 1035 87 1037
rect 193 1039 199 1041
rect 193 1037 195 1039
rect 197 1037 199 1039
rect 193 1020 199 1037
rect 301 1039 307 1041
rect 301 1037 303 1039
rect 305 1037 307 1039
rect 301 1035 307 1037
rect 512 1039 530 1041
rect 512 1037 514 1039
rect 516 1037 526 1039
rect 528 1037 530 1039
rect 512 1035 530 1037
rect 576 1039 582 1041
rect 576 1037 578 1039
rect 580 1037 582 1039
rect 576 1026 582 1037
rect 656 1039 662 1041
rect 656 1037 658 1039
rect 660 1037 662 1039
rect 656 1035 662 1037
rect 674 1039 692 1041
rect 674 1037 676 1039
rect 678 1037 688 1039
rect 690 1037 692 1039
rect 674 1035 692 1037
rect 700 1039 706 1041
rect 700 1037 702 1039
rect 704 1037 706 1039
rect 700 1026 706 1037
rect 101 907 107 909
rect 101 905 103 907
rect 105 905 107 907
rect 101 903 107 905
rect 117 907 135 909
rect 117 905 119 907
rect 121 905 131 907
rect 133 905 135 907
rect 117 903 135 905
rect 145 907 151 909
rect 145 905 147 907
rect 149 905 151 907
rect 145 903 151 905
rect 253 907 259 909
rect 253 905 255 907
rect 257 905 259 907
rect 253 903 259 905
rect 297 907 303 909
rect 297 905 299 907
rect 301 905 303 907
rect 297 903 303 905
rect 564 907 570 909
rect 564 905 566 907
rect 568 905 570 907
rect 564 903 570 905
rect 580 907 586 909
rect 580 905 582 907
rect 584 905 586 907
rect 580 903 586 905
rect 624 907 630 909
rect 624 905 626 907
rect 628 905 630 907
rect 624 903 630 905
rect 736 907 742 909
rect 736 905 738 907
rect 740 905 742 907
rect 736 903 742 905
rect 117 895 123 897
rect 117 893 119 895
rect 121 893 123 895
rect 117 891 123 893
rect 166 895 172 897
rect 166 893 168 895
rect 170 893 172 895
rect 166 891 172 893
rect 247 895 253 897
rect 247 893 249 895
rect 251 893 253 895
rect 247 891 253 893
rect 265 895 283 897
rect 265 893 267 895
rect 269 893 279 895
rect 281 893 283 895
rect 265 891 283 893
rect 293 895 299 897
rect 293 893 295 895
rect 297 893 299 895
rect 293 891 299 893
rect 337 895 343 897
rect 337 893 339 895
rect 341 893 343 895
rect 337 891 343 893
rect 515 895 521 897
rect 515 893 517 895
rect 519 893 521 895
rect 515 891 521 893
rect 532 895 550 897
rect 532 893 534 895
rect 536 893 546 895
rect 548 893 550 895
rect 532 891 550 893
rect 588 895 594 897
rect 588 893 590 895
rect 592 893 594 895
rect 588 891 594 893
rect 608 895 614 897
rect 608 893 610 895
rect 612 893 614 895
rect 608 891 614 893
rect 692 895 698 897
rect 692 893 694 895
rect 696 893 698 895
rect 692 891 698 893
rect 125 763 131 765
rect 125 761 127 763
rect 129 761 131 763
rect 125 759 131 761
rect 209 763 215 765
rect 209 761 211 763
rect 213 761 215 763
rect 209 759 215 761
rect 229 763 235 765
rect 229 761 231 763
rect 233 761 235 763
rect 229 759 235 761
rect 273 763 291 765
rect 273 761 275 763
rect 277 761 287 763
rect 289 761 291 763
rect 273 759 291 761
rect 302 763 308 765
rect 302 761 304 763
rect 306 761 308 763
rect 302 759 308 761
rect 480 763 486 765
rect 480 761 482 763
rect 484 761 486 763
rect 480 759 486 761
rect 524 763 530 765
rect 524 761 526 763
rect 528 761 530 763
rect 524 759 530 761
rect 540 763 558 765
rect 540 761 542 763
rect 544 761 554 763
rect 556 761 558 763
rect 540 759 558 761
rect 570 763 576 765
rect 570 761 572 763
rect 574 761 576 763
rect 570 759 576 761
rect 651 763 657 765
rect 651 761 653 763
rect 655 761 657 763
rect 651 759 657 761
rect 700 763 706 765
rect 700 761 702 763
rect 704 761 706 763
rect 700 759 706 761
rect 81 751 87 753
rect 81 749 83 751
rect 85 749 87 751
rect 81 747 87 749
rect 193 751 199 753
rect 193 749 195 751
rect 197 749 199 751
rect 193 747 199 749
rect 237 751 243 753
rect 237 749 239 751
rect 241 749 243 751
rect 237 747 243 749
rect 253 751 259 753
rect 253 749 255 751
rect 257 749 259 751
rect 253 747 259 749
rect 321 751 339 753
rect 321 749 323 751
rect 325 749 335 751
rect 337 749 339 751
rect 321 747 339 749
rect 520 751 526 753
rect 520 749 522 751
rect 524 749 526 751
rect 520 747 526 749
rect 564 751 570 753
rect 564 749 566 751
rect 568 749 570 751
rect 564 747 570 749
rect 672 751 678 753
rect 672 749 674 751
rect 676 749 678 751
rect 672 747 678 749
rect 688 751 706 753
rect 688 749 690 751
rect 692 749 702 751
rect 704 749 706 751
rect 688 747 706 749
rect 716 751 722 753
rect 716 749 718 751
rect 720 749 722 751
rect 716 747 722 749
rect 117 619 123 630
rect 117 617 119 619
rect 121 617 123 619
rect 117 615 123 617
rect 131 619 149 621
rect 131 617 133 619
rect 135 617 145 619
rect 147 617 149 619
rect 131 615 149 617
rect 161 619 167 621
rect 161 617 163 619
rect 165 617 167 619
rect 161 615 167 617
rect 241 619 247 630
rect 241 617 243 619
rect 245 617 247 619
rect 241 615 247 617
rect 516 619 522 621
rect 516 617 518 619
rect 520 617 522 619
rect 516 615 522 617
rect 624 619 630 636
rect 624 617 626 619
rect 628 617 630 619
rect 624 615 630 617
rect 736 619 742 621
rect 736 617 738 619
rect 740 617 742 619
rect 736 615 742 617
rect 81 607 87 609
rect 81 605 83 607
rect 85 605 87 607
rect 81 603 87 605
rect 215 607 221 609
rect 215 605 217 607
rect 219 605 221 607
rect 215 603 221 605
rect 235 607 253 609
rect 235 605 237 607
rect 239 605 249 607
rect 251 605 253 607
rect 235 603 253 605
rect 496 607 502 609
rect 496 605 498 607
rect 500 605 502 607
rect 496 588 502 605
rect 628 607 634 609
rect 628 605 630 607
rect 632 605 634 607
rect 628 603 634 605
rect 672 607 678 609
rect 672 605 674 607
rect 676 605 678 607
rect 672 603 678 605
rect 688 607 706 609
rect 688 605 690 607
rect 692 605 702 607
rect 704 605 706 607
rect 688 603 706 605
rect 117 475 123 486
rect 117 473 119 475
rect 121 473 123 475
rect 117 471 123 473
rect 129 475 147 477
rect 129 473 131 475
rect 133 473 143 475
rect 145 473 147 475
rect 129 471 147 473
rect 212 475 218 477
rect 212 473 214 475
rect 216 473 218 475
rect 212 471 218 473
rect 230 475 256 477
rect 230 473 232 475
rect 234 473 252 475
rect 254 473 256 475
rect 230 471 256 473
rect 446 475 464 477
rect 446 473 448 475
rect 450 473 460 475
rect 462 473 464 475
rect 446 471 464 473
rect 588 475 594 477
rect 588 473 590 475
rect 592 473 594 475
rect 588 471 594 473
rect 632 475 638 477
rect 632 473 634 475
rect 636 473 638 475
rect 632 471 638 473
rect 648 475 654 477
rect 648 473 650 475
rect 652 473 654 475
rect 648 471 654 473
rect 736 475 742 477
rect 736 473 738 475
rect 740 473 742 475
rect 736 471 742 473
rect 6 360 19 362
rect 6 358 8 360
rect 10 358 15 360
rect 17 358 19 360
rect 6 356 19 358
rect 106 360 119 362
rect 106 358 108 360
rect 110 358 115 360
rect 117 358 119 360
rect 106 356 119 358
rect 206 360 219 362
rect 206 358 208 360
rect 210 358 215 360
rect 217 358 219 360
rect 206 356 219 358
rect 306 360 319 362
rect 306 358 308 360
rect 310 358 315 360
rect 317 358 319 360
rect 306 356 319 358
rect 406 360 419 362
rect 406 358 408 360
rect 410 358 415 360
rect 417 358 419 360
rect 406 356 419 358
rect 506 360 519 362
rect 506 358 508 360
rect 510 358 515 360
rect 517 358 519 360
rect 506 356 519 358
rect 606 360 619 362
rect 606 358 608 360
rect 610 358 615 360
rect 617 358 619 360
rect 606 356 619 358
rect 706 360 719 362
rect 706 358 708 360
rect 710 358 715 360
rect 717 358 719 360
rect 706 356 719 358
rect 83 228 96 230
rect 83 226 85 228
rect 87 226 92 228
rect 94 226 96 228
rect 83 224 96 226
rect 183 228 196 230
rect 183 226 185 228
rect 187 226 192 228
rect 194 226 196 228
rect 183 224 196 226
rect 283 228 296 230
rect 283 226 285 228
rect 287 226 292 228
rect 294 226 296 228
rect 283 224 296 226
rect 383 228 396 230
rect 383 226 385 228
rect 387 226 392 228
rect 394 226 396 228
rect 383 224 396 226
rect 485 228 498 230
rect 485 226 487 228
rect 489 226 494 228
rect 496 226 498 228
rect 485 224 498 226
rect 585 228 598 230
rect 585 226 587 228
rect 589 226 594 228
rect 596 226 598 228
rect 585 224 598 226
rect 685 228 698 230
rect 685 226 687 228
rect 689 226 694 228
rect 696 226 698 228
rect 685 224 698 226
rect 785 228 798 230
rect 785 226 787 228
rect 789 226 794 228
rect 796 226 798 228
rect 785 224 798 226
rect 83 216 96 218
rect 83 214 85 216
rect 87 214 92 216
rect 94 214 96 216
rect 83 212 96 214
rect 183 216 196 218
rect 183 214 185 216
rect 187 214 192 216
rect 194 214 196 216
rect 183 212 196 214
rect 283 216 296 218
rect 283 214 285 216
rect 287 214 292 216
rect 294 214 296 216
rect 283 212 296 214
rect 383 216 396 218
rect 383 214 385 216
rect 387 214 392 216
rect 394 214 396 216
rect 383 212 396 214
rect 485 216 498 218
rect 485 214 487 216
rect 489 214 494 216
rect 496 214 498 216
rect 485 212 498 214
rect 585 216 598 218
rect 585 214 587 216
rect 589 214 594 216
rect 596 214 598 216
rect 585 212 598 214
rect 685 216 698 218
rect 685 214 687 216
rect 689 214 694 216
rect 696 214 698 216
rect 685 212 698 214
rect 785 216 798 218
rect 785 214 787 216
rect 789 214 794 216
rect 796 214 798 216
rect 785 212 798 214
rect 83 84 96 86
rect 83 82 85 84
rect 87 82 92 84
rect 94 82 96 84
rect 83 80 96 82
rect 183 84 196 86
rect 183 82 185 84
rect 187 82 192 84
rect 194 82 196 84
rect 183 80 196 82
rect 283 84 296 86
rect 283 82 285 84
rect 287 82 292 84
rect 294 82 296 84
rect 283 80 296 82
rect 383 84 396 86
rect 383 82 385 84
rect 387 82 392 84
rect 394 82 396 84
rect 383 80 396 82
rect 485 84 498 86
rect 485 82 487 84
rect 489 82 494 84
rect 496 82 498 84
rect 485 80 498 82
rect 585 84 598 86
rect 585 82 587 84
rect 589 82 594 84
rect 596 82 598 84
rect 585 80 598 82
rect 685 84 698 86
rect 685 82 687 84
rect 689 82 694 84
rect 696 82 698 84
rect 685 80 698 82
rect 785 84 798 86
rect 785 82 787 84
rect 789 82 794 84
rect 796 82 798 84
rect 785 80 798 82
rect 6 72 19 74
rect 6 70 8 72
rect 10 70 15 72
rect 17 70 19 72
rect 6 68 19 70
rect 106 72 119 74
rect 106 70 108 72
rect 110 70 115 72
rect 117 70 119 72
rect 106 68 119 70
rect 206 72 219 74
rect 206 70 208 72
rect 210 70 215 72
rect 217 70 219 72
rect 206 68 219 70
rect 306 72 319 74
rect 306 70 308 72
rect 310 70 315 72
rect 317 70 319 72
rect 306 68 319 70
rect 406 72 419 74
rect 406 70 408 72
rect 410 70 415 72
rect 417 70 419 72
rect 406 68 419 70
rect 506 72 519 74
rect 506 70 508 72
rect 510 70 515 72
rect 517 70 519 72
rect 506 68 519 70
rect 606 72 619 74
rect 606 70 608 72
rect 610 70 615 72
rect 617 70 619 72
rect 606 68 619 70
rect 706 72 719 74
rect 706 70 708 72
rect 710 70 715 72
rect 717 70 719 72
rect 706 68 719 70
rect -11 -88 2 -86
rect -11 -90 -9 -88
rect -7 -90 -2 -88
rect 0 -90 2 -88
rect -11 -92 2 -90
rect 95 -88 108 -86
rect 95 -90 97 -88
rect 99 -90 104 -88
rect 106 -90 108 -88
rect 95 -92 108 -90
rect 201 -88 214 -86
rect 201 -90 203 -88
rect 205 -90 210 -88
rect 212 -90 214 -88
rect 201 -92 214 -90
rect 307 -88 320 -86
rect 307 -90 309 -88
rect 311 -90 316 -88
rect 318 -90 320 -88
rect 307 -92 320 -90
rect 413 -88 426 -86
rect 413 -90 415 -88
rect 417 -90 422 -88
rect 424 -90 426 -88
rect 413 -92 426 -90
rect 519 -88 532 -86
rect 519 -90 521 -88
rect 523 -90 528 -88
rect 530 -90 532 -88
rect 519 -92 532 -90
rect 625 -88 638 -86
rect 625 -90 627 -88
rect 629 -90 634 -88
rect 636 -90 638 -88
rect 625 -92 638 -90
rect 731 -88 744 -86
rect 731 -90 733 -88
rect 735 -90 740 -88
rect 742 -90 744 -88
rect 731 -92 744 -90
rect 837 -88 850 -86
rect 837 -90 839 -88
rect 841 -90 846 -88
rect 848 -90 850 -88
rect 837 -92 850 -90
<< ntie >>
rect 114 1123 120 1125
rect 114 1121 116 1123
rect 118 1121 120 1123
rect 185 1123 191 1125
rect 114 1119 120 1121
rect 185 1121 187 1123
rect 189 1121 191 1123
rect 262 1123 268 1125
rect 185 1119 191 1121
rect 262 1121 264 1123
rect 266 1121 268 1123
rect 262 1119 268 1121
rect 359 1123 377 1125
rect 586 1123 592 1125
rect 359 1121 361 1123
rect 363 1121 373 1123
rect 375 1121 377 1123
rect 359 1119 377 1121
rect 586 1121 588 1123
rect 590 1121 592 1123
rect 638 1123 644 1125
rect 586 1119 592 1121
rect 638 1121 640 1123
rect 642 1121 644 1123
rect 676 1123 694 1125
rect 638 1119 644 1121
rect 676 1121 678 1123
rect 680 1121 690 1123
rect 692 1121 694 1123
rect 676 1119 694 1121
rect 117 1111 135 1113
rect 117 1109 119 1111
rect 121 1109 131 1111
rect 133 1109 135 1111
rect 117 1107 135 1109
rect 145 1111 151 1113
rect 145 1109 147 1111
rect 149 1109 151 1111
rect 145 1107 151 1109
rect 233 1111 239 1113
rect 233 1109 235 1111
rect 237 1109 239 1111
rect 233 1107 239 1109
rect 299 1111 327 1113
rect 299 1109 301 1111
rect 303 1109 323 1111
rect 325 1109 327 1111
rect 299 1107 327 1109
rect 570 1111 588 1113
rect 570 1109 572 1111
rect 574 1109 584 1111
rect 586 1109 588 1111
rect 570 1107 588 1109
rect 602 1111 608 1113
rect 602 1109 604 1111
rect 606 1109 608 1111
rect 703 1111 709 1113
rect 602 1107 608 1109
rect 703 1109 705 1111
rect 707 1109 709 1111
rect 703 1107 709 1109
rect 114 979 120 981
rect 114 977 116 979
rect 118 977 120 979
rect 257 979 263 981
rect 114 975 120 977
rect 257 977 259 979
rect 261 977 263 979
rect 257 975 263 977
rect 512 979 530 981
rect 512 977 514 979
rect 516 977 526 979
rect 528 977 530 979
rect 656 979 662 981
rect 512 975 530 977
rect 656 977 658 979
rect 660 977 662 979
rect 656 975 662 977
rect 674 979 692 981
rect 674 977 676 979
rect 678 977 688 979
rect 690 977 692 979
rect 674 975 692 977
rect 117 967 135 969
rect 117 965 119 967
rect 121 965 131 967
rect 133 965 135 967
rect 117 963 135 965
rect 145 967 151 969
rect 145 965 147 967
rect 149 965 151 967
rect 220 967 226 969
rect 145 963 151 965
rect 220 965 222 967
rect 224 965 226 967
rect 297 967 303 969
rect 220 963 226 965
rect 297 965 299 967
rect 301 965 303 967
rect 531 967 537 969
rect 297 963 303 965
rect 531 965 533 967
rect 535 965 537 967
rect 580 967 586 969
rect 531 963 537 965
rect 580 965 582 967
rect 584 965 586 967
rect 580 963 586 965
rect 624 967 638 969
rect 624 965 626 967
rect 628 965 634 967
rect 636 965 638 967
rect 703 967 709 969
rect 624 963 638 965
rect 703 965 705 967
rect 707 965 709 967
rect 703 963 709 965
rect 82 835 96 837
rect 82 833 84 835
rect 86 833 92 835
rect 94 833 96 835
rect 82 831 96 833
rect 117 835 123 837
rect 117 833 119 835
rect 121 833 123 835
rect 117 831 123 833
rect 166 835 172 837
rect 166 833 168 835
rect 170 833 172 835
rect 166 831 172 833
rect 247 835 253 837
rect 247 833 249 835
rect 251 833 253 835
rect 247 831 253 833
rect 265 835 283 837
rect 265 833 267 835
rect 269 833 279 835
rect 281 833 283 835
rect 265 831 283 833
rect 293 835 299 837
rect 293 833 295 835
rect 297 833 299 835
rect 293 831 299 833
rect 381 835 387 837
rect 381 833 383 835
rect 385 833 387 835
rect 381 831 387 833
rect 515 835 521 837
rect 515 833 517 835
rect 519 833 521 835
rect 515 831 521 833
rect 532 835 550 837
rect 532 833 534 835
rect 536 833 546 835
rect 548 833 550 835
rect 532 831 550 833
rect 588 835 594 837
rect 588 833 590 835
rect 592 833 594 835
rect 588 831 594 833
rect 608 835 614 837
rect 608 833 610 835
rect 612 833 614 835
rect 608 831 614 833
rect 648 835 654 837
rect 648 833 650 835
rect 652 833 654 835
rect 648 831 654 833
rect 169 823 175 825
rect 169 821 171 823
rect 173 821 175 823
rect 169 819 175 821
rect 209 823 215 825
rect 209 821 211 823
rect 213 821 215 823
rect 209 819 215 821
rect 229 823 235 825
rect 229 821 231 823
rect 233 821 235 823
rect 229 819 235 821
rect 273 823 291 825
rect 273 821 275 823
rect 277 821 287 823
rect 289 821 291 823
rect 273 819 291 821
rect 302 823 308 825
rect 302 821 304 823
rect 306 821 308 823
rect 302 819 308 821
rect 436 823 442 825
rect 436 821 438 823
rect 440 821 442 823
rect 436 819 442 821
rect 524 823 530 825
rect 524 821 526 823
rect 528 821 530 823
rect 524 819 530 821
rect 540 823 558 825
rect 540 821 542 823
rect 544 821 554 823
rect 556 821 558 823
rect 540 819 558 821
rect 570 823 576 825
rect 570 821 572 823
rect 574 821 576 823
rect 570 819 576 821
rect 651 823 657 825
rect 651 821 653 823
rect 655 821 657 823
rect 651 819 657 821
rect 700 823 706 825
rect 700 821 702 823
rect 704 821 706 823
rect 700 819 706 821
rect 727 823 741 825
rect 727 821 729 823
rect 731 821 737 823
rect 739 821 741 823
rect 727 819 741 821
rect 114 691 120 693
rect 114 689 116 691
rect 118 689 120 691
rect 185 691 199 693
rect 114 687 120 689
rect 185 689 187 691
rect 189 689 195 691
rect 197 689 199 691
rect 185 687 199 689
rect 237 691 243 693
rect 237 689 239 691
rect 241 689 243 691
rect 286 691 292 693
rect 237 687 243 689
rect 286 689 288 691
rect 290 689 292 691
rect 321 691 339 693
rect 286 687 292 689
rect 321 689 323 691
rect 325 689 335 691
rect 337 689 339 691
rect 321 687 339 689
rect 520 691 526 693
rect 520 689 522 691
rect 524 689 526 691
rect 597 691 603 693
rect 520 687 526 689
rect 597 689 599 691
rect 601 689 603 691
rect 672 691 678 693
rect 597 687 603 689
rect 672 689 674 691
rect 676 689 678 691
rect 672 687 678 689
rect 688 691 706 693
rect 688 689 690 691
rect 692 689 702 691
rect 704 689 706 691
rect 688 687 706 689
rect 131 679 149 681
rect 131 677 133 679
rect 135 677 145 679
rect 147 677 149 679
rect 131 675 149 677
rect 161 679 167 681
rect 161 677 163 679
rect 165 677 167 679
rect 161 675 167 677
rect 560 679 566 681
rect 560 677 562 679
rect 564 677 566 679
rect 703 679 709 681
rect 560 675 566 677
rect 703 677 705 679
rect 707 677 709 679
rect 703 675 709 677
rect 114 547 120 549
rect 114 545 116 547
rect 118 545 120 547
rect 215 547 221 549
rect 114 543 120 545
rect 215 545 217 547
rect 219 545 221 547
rect 215 543 221 545
rect 235 547 253 549
rect 235 545 237 547
rect 239 545 249 547
rect 251 545 253 547
rect 235 543 253 545
rect 496 547 524 549
rect 496 545 498 547
rect 500 545 520 547
rect 522 545 524 547
rect 496 543 524 545
rect 584 547 590 549
rect 584 545 586 547
rect 588 545 590 547
rect 584 543 590 545
rect 672 547 678 549
rect 672 545 674 547
rect 676 545 678 547
rect 672 543 678 545
rect 688 547 706 549
rect 688 545 690 547
rect 692 545 702 547
rect 704 545 706 547
rect 688 543 706 545
rect 129 535 147 537
rect 129 533 131 535
rect 133 533 143 535
rect 145 533 147 535
rect 179 535 185 537
rect 129 531 147 533
rect 179 533 181 535
rect 183 533 185 535
rect 231 535 237 537
rect 179 531 185 533
rect 231 533 233 535
rect 235 533 237 535
rect 446 535 464 537
rect 446 533 448 535
rect 450 533 460 535
rect 462 533 464 535
rect 231 531 237 533
rect 446 531 464 533
rect 555 535 561 537
rect 555 533 557 535
rect 559 533 561 535
rect 632 535 638 537
rect 555 531 561 533
rect 632 533 634 535
rect 636 533 638 535
rect 703 535 709 537
rect 632 531 638 533
rect 703 533 705 535
rect 707 533 709 535
rect 703 531 709 533
rect 6 300 12 302
rect 6 298 8 300
rect 10 298 12 300
rect 6 296 12 298
rect 106 300 112 302
rect 106 298 108 300
rect 110 298 112 300
rect 106 296 112 298
rect 206 300 212 302
rect 206 298 208 300
rect 210 298 212 300
rect 206 296 212 298
rect 306 300 312 302
rect 306 298 308 300
rect 310 298 312 300
rect 306 296 312 298
rect 406 300 412 302
rect 406 298 408 300
rect 410 298 412 300
rect 406 296 412 298
rect 506 300 512 302
rect 506 298 508 300
rect 510 298 512 300
rect 506 296 512 298
rect 606 300 612 302
rect 606 298 608 300
rect 610 298 612 300
rect 606 296 612 298
rect 706 300 712 302
rect 706 298 708 300
rect 710 298 712 300
rect 706 296 712 298
rect 90 288 96 290
rect 90 286 92 288
rect 94 286 96 288
rect 90 284 96 286
rect 190 288 196 290
rect 190 286 192 288
rect 194 286 196 288
rect 190 284 196 286
rect 290 288 296 290
rect 290 286 292 288
rect 294 286 296 288
rect 290 284 296 286
rect 390 288 396 290
rect 390 286 392 288
rect 394 286 396 288
rect 390 284 396 286
rect 492 288 498 290
rect 492 286 494 288
rect 496 286 498 288
rect 492 284 498 286
rect 592 288 598 290
rect 592 286 594 288
rect 596 286 598 288
rect 592 284 598 286
rect 692 288 698 290
rect 692 286 694 288
rect 696 286 698 288
rect 692 284 698 286
rect 792 288 798 290
rect 792 286 794 288
rect 796 286 798 288
rect 792 284 798 286
rect 90 156 96 158
rect 90 154 92 156
rect 94 154 96 156
rect 90 152 96 154
rect 190 156 196 158
rect 190 154 192 156
rect 194 154 196 156
rect 190 152 196 154
rect 290 156 296 158
rect 290 154 292 156
rect 294 154 296 156
rect 290 152 296 154
rect 390 156 396 158
rect 390 154 392 156
rect 394 154 396 156
rect 390 152 396 154
rect 492 156 498 158
rect 492 154 494 156
rect 496 154 498 156
rect 492 152 498 154
rect 592 156 598 158
rect 592 154 594 156
rect 596 154 598 156
rect 592 152 598 154
rect 692 156 698 158
rect 692 154 694 156
rect 696 154 698 156
rect 692 152 698 154
rect 792 156 798 158
rect 792 154 794 156
rect 796 154 798 156
rect 792 152 798 154
rect 90 144 96 146
rect 90 142 92 144
rect 94 142 96 144
rect 90 140 96 142
rect 190 144 196 146
rect 190 142 192 144
rect 194 142 196 144
rect 190 140 196 142
rect 290 144 296 146
rect 290 142 292 144
rect 294 142 296 144
rect 290 140 296 142
rect 390 144 396 146
rect 390 142 392 144
rect 394 142 396 144
rect 390 140 396 142
rect 492 144 498 146
rect 492 142 494 144
rect 496 142 498 144
rect 492 140 498 142
rect 592 144 598 146
rect 592 142 594 144
rect 596 142 598 144
rect 592 140 598 142
rect 692 144 698 146
rect 692 142 694 144
rect 696 142 698 144
rect 692 140 698 142
rect 792 144 798 146
rect 792 142 794 144
rect 796 142 798 144
rect 792 140 798 142
rect 6 12 12 14
rect 6 10 8 12
rect 10 10 12 12
rect 6 8 12 10
rect 106 12 112 14
rect 106 10 108 12
rect 110 10 112 12
rect 106 8 112 10
rect 206 12 212 14
rect 206 10 208 12
rect 210 10 212 12
rect 206 8 212 10
rect 306 12 312 14
rect 306 10 308 12
rect 310 10 312 12
rect 306 8 312 10
rect 406 12 412 14
rect 406 10 408 12
rect 410 10 412 12
rect 406 8 412 10
rect 506 12 512 14
rect 506 10 508 12
rect 510 10 512 12
rect 506 8 512 10
rect 606 12 612 14
rect 606 10 608 12
rect 610 10 612 12
rect 606 8 612 10
rect 706 12 712 14
rect 706 10 708 12
rect 710 10 712 12
rect 706 8 712 10
rect -11 -28 -5 -26
rect -11 -30 -9 -28
rect -7 -30 -5 -28
rect -11 -32 -5 -30
rect 95 -28 101 -26
rect 95 -30 97 -28
rect 99 -30 101 -28
rect 95 -32 101 -30
rect 201 -28 207 -26
rect 201 -30 203 -28
rect 205 -30 207 -28
rect 201 -32 207 -30
rect 307 -28 313 -26
rect 307 -30 309 -28
rect 311 -30 313 -28
rect 307 -32 313 -30
rect 413 -28 419 -26
rect 413 -30 415 -28
rect 417 -30 419 -28
rect 413 -32 419 -30
rect 519 -28 525 -26
rect 519 -30 521 -28
rect 523 -30 525 -28
rect 519 -32 525 -30
rect 625 -28 631 -26
rect 625 -30 627 -28
rect 629 -30 631 -28
rect 625 -32 631 -30
rect 731 -28 737 -26
rect 731 -30 733 -28
rect 735 -30 737 -28
rect 731 -32 737 -30
rect 837 -28 843 -26
rect 837 -30 839 -28
rect 841 -30 843 -28
rect 837 -32 843 -30
<< nmos >>
rect 87 1162 89 1171
rect 103 1167 105 1176
rect 113 1167 115 1176
rect 123 1167 125 1179
rect 130 1167 132 1179
rect 156 1168 158 1176
rect 167 1165 169 1173
rect 191 1164 193 1173
rect 204 1164 206 1175
rect 211 1164 213 1175
rect 235 1162 237 1171
rect 251 1167 253 1176
rect 261 1167 263 1176
rect 271 1167 273 1179
rect 278 1167 280 1179
rect 311 1162 313 1182
rect 318 1162 320 1182
rect 325 1162 327 1182
rect 332 1162 334 1182
rect 365 1162 367 1171
rect 574 1162 576 1172
rect 584 1162 586 1172
rect 611 1162 613 1171
rect 627 1167 629 1176
rect 637 1167 639 1176
rect 647 1167 649 1179
rect 654 1167 656 1179
rect 682 1162 684 1171
rect 722 1167 724 1182
rect 732 1167 734 1182
rect 90 1050 92 1070
rect 97 1050 99 1070
rect 123 1061 125 1070
rect 151 1059 153 1068
rect 164 1057 166 1068
rect 171 1057 173 1068
rect 195 1060 197 1069
rect 208 1056 210 1069
rect 215 1056 217 1069
rect 222 1056 224 1069
rect 263 1056 265 1062
rect 273 1056 275 1062
rect 285 1056 287 1062
rect 295 1056 297 1062
rect 580 1061 582 1070
rect 608 1059 610 1068
rect 621 1057 623 1068
rect 628 1057 630 1068
rect 656 1050 658 1070
rect 663 1050 665 1070
rect 691 1053 693 1065
rect 698 1053 700 1065
rect 708 1056 710 1065
rect 718 1056 720 1065
rect 734 1061 736 1070
rect 87 1018 89 1027
rect 103 1023 105 1032
rect 113 1023 115 1032
rect 123 1023 125 1035
rect 130 1023 132 1035
rect 158 1018 160 1038
rect 165 1018 167 1038
rect 217 1026 219 1036
rect 227 1026 229 1036
rect 239 1026 241 1036
rect 272 1019 274 1032
rect 279 1019 281 1032
rect 286 1019 288 1032
rect 299 1019 301 1028
rect 518 1018 520 1027
rect 598 1023 600 1038
rect 608 1023 610 1038
rect 634 1020 636 1031
rect 641 1020 643 1031
rect 654 1020 656 1029
rect 680 1018 682 1027
rect 722 1023 724 1038
rect 732 1023 734 1038
rect 88 912 90 920
rect 99 915 101 923
rect 123 917 125 926
rect 151 915 153 924
rect 164 913 166 924
rect 171 913 173 924
rect 208 909 210 921
rect 215 909 217 921
rect 225 912 227 921
rect 235 912 237 921
rect 251 917 253 926
rect 275 913 277 924
rect 282 913 284 924
rect 295 915 297 924
rect 519 909 521 921
rect 526 909 528 921
rect 536 912 538 921
rect 546 912 548 921
rect 562 917 564 926
rect 586 915 588 924
rect 599 913 601 924
rect 606 913 608 924
rect 630 915 632 926
rect 641 907 643 926
rect 651 911 653 926
rect 661 911 663 926
rect 691 909 693 921
rect 698 909 700 921
rect 708 912 710 921
rect 718 912 720 921
rect 734 917 736 926
rect 93 881 95 893
rect 100 881 102 893
rect 123 876 125 885
rect 136 876 138 887
rect 143 876 145 887
rect 172 876 174 885
rect 185 876 187 887
rect 192 876 194 887
rect 225 876 227 887
rect 232 876 234 887
rect 245 876 247 885
rect 271 874 273 883
rect 299 876 301 885
rect 312 876 314 887
rect 319 876 321 887
rect 343 875 345 884
rect 356 875 358 888
rect 363 875 365 888
rect 370 875 372 888
rect 493 876 495 887
rect 500 876 502 887
rect 513 876 515 885
rect 538 874 540 883
rect 566 876 568 887
rect 573 876 575 887
rect 586 876 588 885
rect 614 876 616 885
rect 627 876 629 887
rect 634 876 636 887
rect 663 875 665 888
rect 670 875 672 888
rect 677 875 679 888
rect 690 875 692 884
rect 717 874 719 894
rect 724 874 726 894
rect 731 874 733 894
rect 90 762 92 782
rect 97 762 99 782
rect 104 762 106 782
rect 131 772 133 781
rect 144 768 146 781
rect 151 768 153 781
rect 158 768 160 781
rect 187 769 189 780
rect 194 769 196 780
rect 207 771 209 780
rect 235 771 237 780
rect 248 769 250 780
rect 255 769 257 780
rect 283 773 285 782
rect 308 771 310 780
rect 321 769 323 780
rect 328 769 330 780
rect 451 768 453 781
rect 458 768 460 781
rect 465 768 467 781
rect 478 772 480 781
rect 502 769 504 780
rect 509 769 511 780
rect 522 771 524 780
rect 550 773 552 782
rect 576 771 578 780
rect 589 769 591 780
rect 596 769 598 780
rect 629 769 631 780
rect 636 769 638 780
rect 649 771 651 780
rect 678 769 680 780
rect 685 769 687 780
rect 698 771 700 780
rect 721 763 723 775
rect 728 763 730 775
rect 87 730 89 739
rect 103 735 105 744
rect 113 735 115 744
rect 123 735 125 747
rect 130 735 132 747
rect 160 730 162 745
rect 170 730 172 745
rect 180 730 182 749
rect 191 730 193 741
rect 215 732 217 743
rect 222 732 224 743
rect 235 732 237 741
rect 259 730 261 739
rect 275 735 277 744
rect 285 735 287 744
rect 295 735 297 747
rect 302 735 304 747
rect 327 730 329 739
rect 526 732 528 741
rect 539 732 541 743
rect 546 732 548 743
rect 570 730 572 739
rect 586 735 588 744
rect 596 735 598 744
rect 606 735 608 747
rect 613 735 615 747
rect 650 732 652 743
rect 657 732 659 743
rect 670 732 672 741
rect 698 730 700 739
rect 722 733 724 741
rect 733 736 735 744
rect 89 618 91 633
rect 99 618 101 633
rect 141 629 143 638
rect 167 627 169 636
rect 180 625 182 636
rect 187 625 189 636
rect 213 618 215 633
rect 223 618 225 633
rect 522 628 524 637
rect 535 624 537 637
rect 542 624 544 637
rect 549 624 551 637
rect 582 620 584 630
rect 594 620 596 630
rect 604 620 606 630
rect 656 618 658 638
rect 663 618 665 638
rect 691 621 693 633
rect 698 621 700 633
rect 708 624 710 633
rect 718 624 720 633
rect 734 629 736 638
rect 87 586 89 595
rect 103 591 105 600
rect 113 591 115 600
rect 123 591 125 603
rect 130 591 132 603
rect 158 586 160 606
rect 165 586 167 606
rect 193 588 195 599
rect 200 588 202 599
rect 213 588 215 597
rect 241 586 243 595
rect 526 594 528 600
rect 536 594 538 600
rect 548 594 550 600
rect 558 594 560 600
rect 599 587 601 600
rect 606 587 608 600
rect 613 587 615 600
rect 626 587 628 596
rect 650 588 652 599
rect 657 588 659 599
rect 670 588 672 597
rect 698 586 700 595
rect 724 586 726 606
rect 731 586 733 606
rect 89 474 91 489
rect 99 474 101 489
rect 139 485 141 494
rect 167 477 169 489
rect 174 477 176 489
rect 184 480 186 489
rect 194 480 196 489
rect 210 485 212 494
rect 237 484 239 494
rect 247 484 249 494
rect 456 485 458 494
rect 489 474 491 494
rect 496 474 498 494
rect 503 474 505 494
rect 510 474 512 494
rect 543 477 545 489
rect 550 477 552 489
rect 560 480 562 489
rect 570 480 572 489
rect 586 485 588 494
rect 610 481 612 492
rect 617 481 619 492
rect 630 483 632 492
rect 654 483 656 491
rect 665 480 667 488
rect 691 477 693 489
rect 698 477 700 489
rect 708 480 710 489
rect 718 480 720 489
rect 734 485 736 494
rect 14 340 16 350
rect 25 340 27 351
rect 35 340 37 351
rect 45 345 47 356
rect 55 342 57 353
rect 75 342 77 352
rect 88 342 90 349
rect 114 340 116 350
rect 125 340 127 351
rect 135 340 137 351
rect 145 345 147 356
rect 155 342 157 353
rect 175 342 177 352
rect 188 342 190 349
rect 214 340 216 350
rect 225 340 227 351
rect 235 340 237 351
rect 245 345 247 356
rect 255 342 257 353
rect 275 342 277 352
rect 288 342 290 349
rect 314 340 316 350
rect 325 340 327 351
rect 335 340 337 351
rect 345 345 347 356
rect 355 342 357 353
rect 375 342 377 352
rect 388 342 390 349
rect 414 340 416 350
rect 425 340 427 351
rect 435 340 437 351
rect 445 345 447 356
rect 455 342 457 353
rect 475 342 477 352
rect 488 342 490 349
rect 514 340 516 350
rect 525 340 527 351
rect 535 340 537 351
rect 545 345 547 356
rect 555 342 557 353
rect 575 342 577 352
rect 588 342 590 349
rect 614 340 616 350
rect 625 340 627 351
rect 635 340 637 351
rect 645 345 647 356
rect 655 342 657 353
rect 675 342 677 352
rect 688 342 690 349
rect 714 340 716 350
rect 725 340 727 351
rect 735 340 737 351
rect 745 345 747 356
rect 755 342 757 353
rect 775 342 777 352
rect 788 342 790 349
rect 12 237 14 244
rect 25 234 27 244
rect 45 233 47 244
rect 55 230 57 241
rect 65 235 67 246
rect 75 235 77 246
rect 86 236 88 246
rect 112 237 114 244
rect 125 234 127 244
rect 145 233 147 244
rect 155 230 157 241
rect 165 235 167 246
rect 175 235 177 246
rect 186 236 188 246
rect 212 237 214 244
rect 225 234 227 244
rect 245 233 247 244
rect 255 230 257 241
rect 265 235 267 246
rect 275 235 277 246
rect 286 236 288 246
rect 312 237 314 244
rect 325 234 327 244
rect 345 233 347 244
rect 355 230 357 241
rect 365 235 367 246
rect 375 235 377 246
rect 386 236 388 246
rect 414 237 416 244
rect 427 234 429 244
rect 447 233 449 244
rect 457 230 459 241
rect 467 235 469 246
rect 477 235 479 246
rect 488 236 490 246
rect 514 237 516 244
rect 527 234 529 244
rect 547 233 549 244
rect 557 230 559 241
rect 567 235 569 246
rect 577 235 579 246
rect 588 236 590 246
rect 614 237 616 244
rect 627 234 629 244
rect 647 233 649 244
rect 657 230 659 241
rect 667 235 669 246
rect 677 235 679 246
rect 688 236 690 246
rect 714 237 716 244
rect 727 234 729 244
rect 747 233 749 244
rect 757 230 759 241
rect 767 235 769 246
rect 777 235 779 246
rect 788 236 790 246
rect 12 198 14 205
rect 25 198 27 208
rect 45 198 47 209
rect 55 201 57 212
rect 65 196 67 207
rect 75 196 77 207
rect 86 196 88 206
rect 112 198 114 205
rect 125 198 127 208
rect 145 198 147 209
rect 155 201 157 212
rect 165 196 167 207
rect 175 196 177 207
rect 186 196 188 206
rect 212 198 214 205
rect 225 198 227 208
rect 245 198 247 209
rect 255 201 257 212
rect 265 196 267 207
rect 275 196 277 207
rect 286 196 288 206
rect 312 198 314 205
rect 325 198 327 208
rect 345 198 347 209
rect 355 201 357 212
rect 365 196 367 207
rect 375 196 377 207
rect 386 196 388 206
rect 414 198 416 205
rect 427 198 429 208
rect 447 198 449 209
rect 457 201 459 212
rect 467 196 469 207
rect 477 196 479 207
rect 488 196 490 206
rect 514 198 516 205
rect 527 198 529 208
rect 547 198 549 209
rect 557 201 559 212
rect 567 196 569 207
rect 577 196 579 207
rect 588 196 590 206
rect 614 198 616 205
rect 627 198 629 208
rect 647 198 649 209
rect 657 201 659 212
rect 667 196 669 207
rect 677 196 679 207
rect 688 196 690 206
rect 714 198 716 205
rect 727 198 729 208
rect 747 198 749 209
rect 757 201 759 212
rect 767 196 769 207
rect 777 196 779 207
rect 788 196 790 206
rect 12 93 14 100
rect 25 90 27 100
rect 45 89 47 100
rect 55 86 57 97
rect 65 91 67 102
rect 75 91 77 102
rect 86 92 88 102
rect 112 93 114 100
rect 125 90 127 100
rect 145 89 147 100
rect 155 86 157 97
rect 165 91 167 102
rect 175 91 177 102
rect 186 92 188 102
rect 212 93 214 100
rect 225 90 227 100
rect 245 89 247 100
rect 255 86 257 97
rect 265 91 267 102
rect 275 91 277 102
rect 286 92 288 102
rect 312 93 314 100
rect 325 90 327 100
rect 345 89 347 100
rect 355 86 357 97
rect 365 91 367 102
rect 375 91 377 102
rect 386 92 388 102
rect 414 93 416 100
rect 427 90 429 100
rect 447 89 449 100
rect 457 86 459 97
rect 467 91 469 102
rect 477 91 479 102
rect 488 92 490 102
rect 514 93 516 100
rect 527 90 529 100
rect 547 89 549 100
rect 557 86 559 97
rect 567 91 569 102
rect 577 91 579 102
rect 588 92 590 102
rect 614 93 616 100
rect 627 90 629 100
rect 647 89 649 100
rect 657 86 659 97
rect 667 91 669 102
rect 677 91 679 102
rect 688 92 690 102
rect 714 93 716 100
rect 727 90 729 100
rect 747 89 749 100
rect 757 86 759 97
rect 767 91 769 102
rect 777 91 779 102
rect 788 92 790 102
rect 14 52 16 62
rect 25 52 27 63
rect 35 52 37 63
rect 45 57 47 68
rect 55 54 57 65
rect 75 54 77 64
rect 88 54 90 61
rect 114 52 116 62
rect 125 52 127 63
rect 135 52 137 63
rect 145 57 147 68
rect 155 54 157 65
rect 175 54 177 64
rect 188 54 190 61
rect 214 52 216 62
rect 225 52 227 63
rect 235 52 237 63
rect 245 57 247 68
rect 255 54 257 65
rect 275 54 277 64
rect 288 54 290 61
rect 314 52 316 62
rect 325 52 327 63
rect 335 52 337 63
rect 345 57 347 68
rect 355 54 357 65
rect 375 54 377 64
rect 388 54 390 61
rect 414 52 416 62
rect 425 52 427 63
rect 435 52 437 63
rect 445 57 447 68
rect 455 54 457 65
rect 475 54 477 64
rect 488 54 490 61
rect 514 52 516 62
rect 525 52 527 63
rect 535 52 537 63
rect 545 57 547 68
rect 555 54 557 65
rect 575 54 577 64
rect 588 54 590 61
rect 614 52 616 62
rect 625 52 627 63
rect 635 52 637 63
rect 645 57 647 68
rect 655 54 657 65
rect 675 54 677 64
rect 688 54 690 61
rect 714 52 716 62
rect 725 52 727 63
rect 735 52 737 63
rect 745 57 747 68
rect 755 54 757 65
rect 775 54 777 64
rect 788 54 790 61
rect -3 -80 -1 -70
rect 8 -81 10 -70
rect 18 -81 20 -70
rect 28 -86 30 -75
rect 38 -83 40 -72
rect 58 -82 60 -72
rect 71 -79 73 -72
rect 103 -80 105 -70
rect 114 -81 116 -70
rect 124 -81 126 -70
rect 134 -86 136 -75
rect 144 -83 146 -72
rect 164 -82 166 -72
rect 177 -79 179 -72
rect 209 -80 211 -70
rect 220 -81 222 -70
rect 230 -81 232 -70
rect 240 -86 242 -75
rect 250 -83 252 -72
rect 270 -82 272 -72
rect 283 -79 285 -72
rect 315 -80 317 -70
rect 326 -81 328 -70
rect 336 -81 338 -70
rect 346 -86 348 -75
rect 356 -83 358 -72
rect 376 -82 378 -72
rect 389 -79 391 -72
rect 421 -80 423 -70
rect 432 -81 434 -70
rect 442 -81 444 -70
rect 452 -86 454 -75
rect 462 -83 464 -72
rect 482 -82 484 -72
rect 495 -79 497 -72
rect 527 -80 529 -70
rect 538 -81 540 -70
rect 548 -81 550 -70
rect 558 -86 560 -75
rect 568 -83 570 -72
rect 588 -82 590 -72
rect 601 -79 603 -72
rect 633 -80 635 -70
rect 644 -81 646 -70
rect 654 -81 656 -70
rect 664 -86 666 -75
rect 674 -83 676 -72
rect 694 -82 696 -72
rect 707 -79 709 -72
rect 739 -80 741 -70
rect 750 -81 752 -70
rect 760 -81 762 -70
rect 770 -86 772 -75
rect 780 -83 782 -72
rect 800 -82 802 -72
rect 813 -79 815 -72
rect 845 -80 847 -70
rect 856 -81 858 -70
rect 866 -81 868 -70
rect 876 -86 878 -75
rect 886 -83 888 -72
rect 906 -82 908 -72
rect 919 -79 921 -72
<< pmos >>
rect 95 1122 97 1149
rect 111 1131 113 1149
rect 121 1131 123 1149
rect 131 1122 133 1149
rect 158 1122 160 1150
rect 165 1122 167 1150
rect 191 1131 193 1149
rect 201 1129 203 1142
rect 211 1129 213 1142
rect 243 1122 245 1149
rect 259 1131 261 1149
rect 269 1131 271 1149
rect 279 1122 281 1149
rect 305 1126 307 1143
rect 315 1126 317 1143
rect 325 1126 327 1143
rect 335 1126 337 1143
rect 365 1132 367 1150
rect 574 1123 576 1147
rect 584 1131 586 1147
rect 619 1122 621 1149
rect 635 1131 637 1149
rect 645 1131 647 1149
rect 655 1122 657 1149
rect 682 1132 684 1150
rect 710 1122 712 1149
rect 717 1122 719 1149
rect 727 1122 729 1149
rect 734 1122 736 1149
rect 87 1086 89 1110
rect 97 1086 99 1110
rect 123 1082 125 1100
rect 151 1083 153 1101
rect 161 1090 163 1103
rect 171 1090 173 1103
rect 195 1084 197 1102
rect 205 1089 207 1102
rect 215 1089 217 1102
rect 227 1088 229 1101
rect 267 1083 269 1108
rect 274 1083 276 1108
rect 281 1083 283 1108
rect 288 1083 290 1108
rect 298 1083 300 1101
rect 305 1083 307 1101
rect 312 1083 314 1101
rect 319 1083 321 1101
rect 580 1082 582 1100
rect 608 1083 610 1101
rect 618 1090 620 1103
rect 628 1090 630 1103
rect 656 1086 658 1110
rect 666 1086 668 1110
rect 690 1083 692 1110
rect 700 1083 702 1101
rect 710 1083 712 1101
rect 726 1083 728 1110
rect 95 978 97 1005
rect 111 987 113 1005
rect 121 987 123 1005
rect 131 978 133 1005
rect 155 978 157 1002
rect 165 978 167 1002
rect 199 978 201 1006
rect 206 978 208 1006
rect 213 978 215 1006
rect 223 978 225 1006
rect 230 978 232 1006
rect 237 978 239 1006
rect 267 987 269 1000
rect 279 986 281 999
rect 289 986 291 999
rect 299 986 301 1004
rect 518 988 520 1006
rect 586 978 588 1005
rect 593 978 595 1005
rect 603 978 605 1005
rect 610 978 612 1005
rect 634 985 636 998
rect 644 985 646 998
rect 654 987 656 1005
rect 680 988 682 1006
rect 710 978 712 1005
rect 717 978 719 1005
rect 727 978 729 1005
rect 734 978 736 1005
rect 90 938 92 966
rect 97 938 99 966
rect 123 938 125 956
rect 151 939 153 957
rect 161 946 163 959
rect 171 946 173 959
rect 207 939 209 966
rect 217 939 219 957
rect 227 939 229 957
rect 243 939 245 966
rect 275 946 277 959
rect 285 946 287 959
rect 295 939 297 957
rect 518 939 520 966
rect 528 939 530 957
rect 538 939 540 957
rect 554 939 556 966
rect 586 939 588 957
rect 596 946 598 959
rect 606 946 608 959
rect 631 939 633 957
rect 641 939 643 957
rect 651 939 653 957
rect 661 939 663 957
rect 690 939 692 966
rect 700 939 702 957
rect 710 939 712 957
rect 726 939 728 966
rect 89 843 91 857
rect 99 843 101 857
rect 123 843 125 861
rect 133 841 135 854
rect 143 841 145 854
rect 172 843 174 861
rect 182 841 184 854
rect 192 841 194 854
rect 225 841 227 854
rect 235 841 237 854
rect 245 843 247 861
rect 271 844 273 862
rect 299 843 301 861
rect 309 841 311 854
rect 319 841 321 854
rect 343 842 345 860
rect 353 842 355 855
rect 363 842 365 855
rect 375 843 377 856
rect 493 841 495 854
rect 503 841 505 854
rect 513 843 515 861
rect 538 844 540 862
rect 566 841 568 854
rect 576 841 578 854
rect 586 843 588 861
rect 614 843 616 861
rect 624 841 626 854
rect 634 841 636 854
rect 658 843 660 856
rect 670 842 672 855
rect 680 842 682 855
rect 690 842 692 860
rect 714 834 716 854
rect 724 834 726 854
rect 734 834 736 854
rect 87 802 89 822
rect 97 802 99 822
rect 107 802 109 822
rect 131 796 133 814
rect 141 801 143 814
rect 151 801 153 814
rect 163 800 165 813
rect 187 802 189 815
rect 197 802 199 815
rect 207 795 209 813
rect 235 795 237 813
rect 245 802 247 815
rect 255 802 257 815
rect 283 794 285 812
rect 308 795 310 813
rect 318 802 320 815
rect 328 802 330 815
rect 446 800 448 813
rect 458 801 460 814
rect 468 801 470 814
rect 478 796 480 814
rect 502 802 504 815
rect 512 802 514 815
rect 522 795 524 813
rect 550 794 552 812
rect 576 795 578 813
rect 586 802 588 815
rect 596 802 598 815
rect 629 802 631 815
rect 639 802 641 815
rect 649 795 651 813
rect 678 802 680 815
rect 688 802 690 815
rect 698 795 700 813
rect 722 799 724 813
rect 732 799 734 813
rect 95 690 97 717
rect 111 699 113 717
rect 121 699 123 717
rect 131 690 133 717
rect 160 699 162 717
rect 170 699 172 717
rect 180 699 182 717
rect 190 699 192 717
rect 215 697 217 710
rect 225 697 227 710
rect 235 699 237 717
rect 267 690 269 717
rect 283 699 285 717
rect 293 699 295 717
rect 303 690 305 717
rect 327 700 329 718
rect 526 699 528 717
rect 536 697 538 710
rect 546 697 548 710
rect 578 690 580 717
rect 594 699 596 717
rect 604 699 606 717
rect 614 690 616 717
rect 650 697 652 710
rect 660 697 662 710
rect 670 699 672 717
rect 698 700 700 718
rect 724 690 726 718
rect 731 690 733 718
rect 87 651 89 678
rect 94 651 96 678
rect 104 651 106 678
rect 111 651 113 678
rect 141 650 143 668
rect 167 651 169 669
rect 177 658 179 671
rect 187 658 189 671
rect 211 651 213 678
rect 218 651 220 678
rect 228 651 230 678
rect 235 651 237 678
rect 522 652 524 670
rect 532 657 534 670
rect 542 657 544 670
rect 554 656 556 669
rect 584 650 586 678
rect 591 650 593 678
rect 598 650 600 678
rect 608 650 610 678
rect 615 650 617 678
rect 622 650 624 678
rect 656 654 658 678
rect 666 654 668 678
rect 690 651 692 678
rect 700 651 702 669
rect 710 651 712 669
rect 726 651 728 678
rect 95 546 97 573
rect 111 555 113 573
rect 121 555 123 573
rect 131 546 133 573
rect 155 546 157 570
rect 165 546 167 570
rect 193 553 195 566
rect 203 553 205 566
rect 213 555 215 573
rect 241 556 243 574
rect 502 555 504 573
rect 509 555 511 573
rect 516 555 518 573
rect 523 555 525 573
rect 533 548 535 573
rect 540 548 542 573
rect 547 548 549 573
rect 554 548 556 573
rect 594 555 596 568
rect 606 554 608 567
rect 616 554 618 567
rect 626 554 628 572
rect 650 553 652 566
rect 660 553 662 566
rect 670 555 672 573
rect 698 556 700 574
rect 724 546 726 570
rect 734 546 736 570
rect 87 507 89 534
rect 94 507 96 534
rect 104 507 106 534
rect 111 507 113 534
rect 139 506 141 524
rect 166 507 168 534
rect 176 507 178 525
rect 186 507 188 525
rect 202 507 204 534
rect 237 509 239 525
rect 247 509 249 533
rect 456 506 458 524
rect 486 513 488 530
rect 496 513 498 530
rect 506 513 508 530
rect 516 513 518 530
rect 542 507 544 534
rect 552 507 554 525
rect 562 507 564 525
rect 578 507 580 534
rect 610 514 612 527
rect 620 514 622 527
rect 630 507 632 525
rect 656 506 658 534
rect 663 506 665 534
rect 690 507 692 534
rect 700 507 702 525
rect 710 507 712 525
rect 726 507 728 534
rect 12 314 14 327
rect 23 305 25 327
rect 33 305 35 327
rect 43 305 45 327
rect 57 305 59 327
rect 75 314 77 327
rect 88 309 90 319
rect 112 314 114 327
rect 123 305 125 327
rect 133 305 135 327
rect 143 305 145 327
rect 157 305 159 327
rect 175 314 177 327
rect 188 309 190 319
rect 212 314 214 327
rect 223 305 225 327
rect 233 305 235 327
rect 243 305 245 327
rect 257 305 259 327
rect 275 314 277 327
rect 288 309 290 319
rect 312 314 314 327
rect 323 305 325 327
rect 333 305 335 327
rect 343 305 345 327
rect 357 305 359 327
rect 375 314 377 327
rect 388 309 390 319
rect 412 314 414 327
rect 423 305 425 327
rect 433 305 435 327
rect 443 305 445 327
rect 457 305 459 327
rect 475 314 477 327
rect 488 309 490 319
rect 512 314 514 327
rect 523 305 525 327
rect 533 305 535 327
rect 543 305 545 327
rect 557 305 559 327
rect 575 314 577 327
rect 588 309 590 319
rect 612 314 614 327
rect 623 305 625 327
rect 633 305 635 327
rect 643 305 645 327
rect 657 305 659 327
rect 675 314 677 327
rect 688 309 690 319
rect 712 314 714 327
rect 723 305 725 327
rect 733 305 735 327
rect 743 305 745 327
rect 757 305 759 327
rect 775 314 777 327
rect 788 309 790 319
rect 12 267 14 277
rect 25 259 27 272
rect 43 259 45 281
rect 57 259 59 281
rect 67 259 69 281
rect 77 259 79 281
rect 88 259 90 272
rect 112 267 114 277
rect 125 259 127 272
rect 143 259 145 281
rect 157 259 159 281
rect 167 259 169 281
rect 177 259 179 281
rect 188 259 190 272
rect 212 267 214 277
rect 225 259 227 272
rect 243 259 245 281
rect 257 259 259 281
rect 267 259 269 281
rect 277 259 279 281
rect 288 259 290 273
rect 312 267 314 277
rect 325 259 327 272
rect 343 259 345 281
rect 357 259 359 281
rect 367 259 369 281
rect 377 259 379 281
rect 388 259 390 272
rect 414 267 416 277
rect 427 259 429 272
rect 445 259 447 281
rect 459 259 461 281
rect 469 259 471 281
rect 479 259 481 281
rect 490 260 492 273
rect 514 267 516 277
rect 527 259 529 272
rect 545 259 547 281
rect 559 259 561 281
rect 569 259 571 281
rect 579 259 581 281
rect 590 259 592 272
rect 614 267 616 277
rect 627 259 629 272
rect 645 259 647 281
rect 659 259 661 281
rect 669 259 671 281
rect 679 259 681 281
rect 690 260 692 273
rect 714 267 716 277
rect 727 259 729 272
rect 745 259 747 281
rect 759 259 761 281
rect 769 259 771 281
rect 779 259 781 281
rect 790 259 792 272
rect 12 165 14 175
rect 25 170 27 183
rect 43 161 45 183
rect 57 161 59 183
rect 67 161 69 183
rect 77 161 79 183
rect 88 170 90 183
rect 112 165 114 175
rect 125 170 127 183
rect 143 161 145 183
rect 157 161 159 183
rect 167 161 169 183
rect 177 161 179 183
rect 188 170 190 183
rect 212 165 214 175
rect 225 170 227 183
rect 243 161 245 183
rect 257 161 259 183
rect 267 161 269 183
rect 277 161 279 183
rect 288 170 290 183
rect 312 165 314 175
rect 325 170 327 183
rect 343 161 345 183
rect 357 161 359 183
rect 367 161 369 183
rect 377 161 379 183
rect 388 170 390 183
rect 414 165 416 175
rect 427 170 429 183
rect 445 161 447 183
rect 459 161 461 183
rect 469 161 471 183
rect 479 161 481 183
rect 490 170 492 183
rect 514 165 516 175
rect 527 170 529 183
rect 545 161 547 183
rect 559 161 561 183
rect 569 161 571 183
rect 579 161 581 183
rect 590 170 592 183
rect 614 165 616 175
rect 627 170 629 183
rect 645 161 647 183
rect 659 161 661 183
rect 669 161 671 183
rect 679 161 681 183
rect 690 170 692 183
rect 714 165 716 175
rect 727 170 729 183
rect 745 161 747 183
rect 759 161 761 183
rect 769 161 771 183
rect 779 161 781 183
rect 790 170 792 183
rect 12 123 14 133
rect 25 115 27 128
rect 43 115 45 137
rect 57 115 59 137
rect 67 115 69 137
rect 77 115 79 137
rect 88 115 90 128
rect 112 123 114 133
rect 125 115 127 128
rect 143 115 145 137
rect 157 115 159 137
rect 167 115 169 137
rect 177 115 179 137
rect 188 115 190 128
rect 212 123 214 133
rect 225 115 227 128
rect 243 115 245 137
rect 257 115 259 137
rect 267 115 269 137
rect 277 115 279 137
rect 288 115 290 128
rect 312 123 314 133
rect 325 115 327 128
rect 343 115 345 137
rect 357 115 359 137
rect 367 115 369 137
rect 377 115 379 137
rect 388 115 390 128
rect 414 123 416 133
rect 427 115 429 128
rect 445 115 447 137
rect 459 115 461 137
rect 469 115 471 137
rect 479 115 481 137
rect 490 115 492 128
rect 514 123 516 133
rect 527 115 529 128
rect 545 115 547 137
rect 559 115 561 137
rect 569 115 571 137
rect 579 115 581 137
rect 590 115 592 128
rect 614 123 616 133
rect 627 115 629 128
rect 645 115 647 137
rect 659 115 661 137
rect 669 115 671 137
rect 679 115 681 137
rect 690 115 692 128
rect 714 123 716 133
rect 727 115 729 128
rect 745 115 747 137
rect 759 115 761 137
rect 769 115 771 137
rect 779 115 781 137
rect 790 115 792 128
rect 12 26 14 39
rect 23 17 25 39
rect 33 17 35 39
rect 43 17 45 39
rect 57 17 59 39
rect 75 26 77 39
rect 88 21 90 31
rect 112 26 114 39
rect 123 17 125 39
rect 133 17 135 39
rect 143 17 145 39
rect 157 17 159 39
rect 175 26 177 39
rect 188 21 190 31
rect 212 26 214 39
rect 223 17 225 39
rect 233 17 235 39
rect 243 17 245 39
rect 257 17 259 39
rect 275 26 277 39
rect 288 21 290 31
rect 312 26 314 39
rect 323 17 325 39
rect 333 17 335 39
rect 343 17 345 39
rect 357 17 359 39
rect 375 26 377 39
rect 388 21 390 31
rect 412 26 414 39
rect 423 17 425 39
rect 433 17 435 39
rect 443 17 445 39
rect 457 17 459 39
rect 475 26 477 39
rect 488 21 490 31
rect 512 26 514 39
rect 523 17 525 39
rect 533 17 535 39
rect 543 17 545 39
rect 557 17 559 39
rect 575 26 577 39
rect 588 21 590 31
rect 612 26 614 39
rect 623 17 625 39
rect 633 17 635 39
rect 643 17 645 39
rect 657 17 659 39
rect 675 26 677 39
rect 688 21 690 31
rect 712 26 714 39
rect 723 17 725 39
rect 733 17 735 39
rect 743 17 745 39
rect 757 17 759 39
rect 775 26 777 39
rect 788 21 790 31
rect -5 -57 -3 -44
rect 6 -57 8 -35
rect 16 -57 18 -35
rect 26 -57 28 -35
rect 40 -57 42 -35
rect 58 -57 60 -44
rect 71 -49 73 -39
rect 101 -57 103 -44
rect 112 -57 114 -35
rect 122 -57 124 -35
rect 132 -57 134 -35
rect 146 -57 148 -35
rect 164 -57 166 -44
rect 177 -49 179 -39
rect 207 -57 209 -44
rect 218 -57 220 -35
rect 228 -57 230 -35
rect 238 -57 240 -35
rect 252 -57 254 -35
rect 270 -57 272 -44
rect 283 -49 285 -39
rect 313 -57 315 -44
rect 324 -57 326 -35
rect 334 -57 336 -35
rect 344 -57 346 -35
rect 358 -57 360 -35
rect 376 -57 378 -44
rect 389 -49 391 -39
rect 419 -57 421 -44
rect 430 -57 432 -35
rect 440 -57 442 -35
rect 450 -57 452 -35
rect 464 -57 466 -35
rect 482 -57 484 -44
rect 495 -49 497 -39
rect 525 -57 527 -44
rect 536 -57 538 -35
rect 546 -57 548 -35
rect 556 -57 558 -35
rect 570 -57 572 -35
rect 588 -57 590 -44
rect 601 -49 603 -39
rect 631 -57 633 -44
rect 642 -57 644 -35
rect 652 -57 654 -35
rect 662 -57 664 -35
rect 676 -57 678 -35
rect 694 -57 696 -44
rect 707 -49 709 -39
rect 737 -57 739 -44
rect 748 -57 750 -35
rect 758 -57 760 -35
rect 768 -57 770 -35
rect 782 -57 784 -35
rect 800 -57 802 -44
rect 813 -49 815 -39
rect 843 -57 845 -44
rect 854 -57 856 -35
rect 864 -57 866 -35
rect 874 -57 876 -35
rect 888 -57 890 -35
rect 906 -57 908 -44
rect 919 -49 921 -39
<< polyct0 >>
rect 119 1155 121 1157
rect 129 1154 131 1156
rect 193 1155 195 1157
rect 267 1155 269 1157
rect 277 1154 279 1156
rect 643 1155 645 1157
rect 327 1148 329 1150
rect 653 1154 655 1156
rect 153 1075 155 1077
rect 197 1075 199 1077
rect 610 1075 612 1077
rect 692 1076 694 1078
rect 702 1075 704 1077
rect 119 1011 121 1013
rect 129 1010 131 1012
rect 297 1011 299 1013
rect 652 1011 654 1013
rect 153 931 155 933
rect 209 932 211 934
rect 219 931 221 933
rect 293 931 295 933
rect 520 932 522 934
rect 530 931 532 933
rect 588 931 590 933
rect 692 932 694 934
rect 702 931 704 933
rect 125 867 127 869
rect 174 867 176 869
rect 243 867 245 869
rect 301 867 303 869
rect 345 867 347 869
rect 511 867 513 869
rect 584 867 586 869
rect 616 867 618 869
rect 688 867 690 869
rect 133 787 135 789
rect 205 787 207 789
rect 237 787 239 789
rect 310 787 312 789
rect 476 787 478 789
rect 520 787 522 789
rect 578 787 580 789
rect 647 787 649 789
rect 696 787 698 789
rect 119 723 121 725
rect 129 722 131 724
rect 233 723 235 725
rect 291 723 293 725
rect 301 722 303 724
rect 528 723 530 725
rect 602 723 604 725
rect 612 722 614 724
rect 668 723 670 725
rect 169 643 171 645
rect 524 643 526 645
rect 692 644 694 646
rect 702 643 704 645
rect 119 579 121 581
rect 129 578 131 580
rect 211 579 213 581
rect 624 579 626 581
rect 668 579 670 581
rect 168 500 170 502
rect 494 506 496 508
rect 178 499 180 501
rect 544 500 546 502
rect 554 499 556 501
rect 628 499 630 501
rect 692 500 694 502
rect 702 499 704 501
rect 23 332 25 334
rect 45 332 47 334
rect 60 332 62 334
rect 123 332 125 334
rect 145 332 147 334
rect 160 332 162 334
rect 223 332 225 334
rect 245 332 247 334
rect 260 332 262 334
rect 323 332 325 334
rect 345 332 347 334
rect 360 332 362 334
rect 423 332 425 334
rect 445 332 447 334
rect 460 332 462 334
rect 523 332 525 334
rect 545 332 547 334
rect 560 332 562 334
rect 623 332 625 334
rect 645 332 647 334
rect 660 332 662 334
rect 723 332 725 334
rect 745 332 747 334
rect 760 332 762 334
rect 40 252 42 254
rect 55 252 57 254
rect 77 252 79 254
rect 140 252 142 254
rect 155 252 157 254
rect 177 252 179 254
rect 240 252 242 254
rect 255 252 257 254
rect 277 252 279 254
rect 340 252 342 254
rect 355 252 357 254
rect 377 252 379 254
rect 442 252 444 254
rect 457 252 459 254
rect 479 252 481 254
rect 542 252 544 254
rect 557 252 559 254
rect 579 252 581 254
rect 642 252 644 254
rect 657 252 659 254
rect 679 252 681 254
rect 742 252 744 254
rect 757 252 759 254
rect 779 252 781 254
rect 40 188 42 190
rect 55 188 57 190
rect 77 188 79 190
rect 140 188 142 190
rect 155 188 157 190
rect 177 188 179 190
rect 240 188 242 190
rect 255 188 257 190
rect 277 188 279 190
rect 340 188 342 190
rect 355 188 357 190
rect 377 188 379 190
rect 442 188 444 190
rect 457 188 459 190
rect 479 188 481 190
rect 542 188 544 190
rect 557 188 559 190
rect 579 188 581 190
rect 642 188 644 190
rect 657 188 659 190
rect 679 188 681 190
rect 742 188 744 190
rect 757 188 759 190
rect 779 188 781 190
rect 40 108 42 110
rect 55 108 57 110
rect 77 108 79 110
rect 140 108 142 110
rect 155 108 157 110
rect 177 108 179 110
rect 240 108 242 110
rect 255 108 257 110
rect 277 108 279 110
rect 340 108 342 110
rect 355 108 357 110
rect 377 108 379 110
rect 442 108 444 110
rect 457 108 459 110
rect 479 108 481 110
rect 542 108 544 110
rect 557 108 559 110
rect 579 108 581 110
rect 642 108 644 110
rect 657 108 659 110
rect 679 108 681 110
rect 742 108 744 110
rect 757 108 759 110
rect 779 108 781 110
rect 23 44 25 46
rect 45 44 47 46
rect 60 44 62 46
rect 123 44 125 46
rect 145 44 147 46
rect 160 44 162 46
rect 223 44 225 46
rect 245 44 247 46
rect 260 44 262 46
rect 323 44 325 46
rect 345 44 347 46
rect 360 44 362 46
rect 423 44 425 46
rect 445 44 447 46
rect 460 44 462 46
rect 523 44 525 46
rect 545 44 547 46
rect 560 44 562 46
rect 623 44 625 46
rect 645 44 647 46
rect 660 44 662 46
rect 723 44 725 46
rect 745 44 747 46
rect 760 44 762 46
rect 6 -64 8 -62
rect 28 -64 30 -62
rect 43 -64 45 -62
rect 112 -64 114 -62
rect 134 -64 136 -62
rect 149 -64 151 -62
rect 218 -64 220 -62
rect 240 -64 242 -62
rect 255 -64 257 -62
rect 324 -64 326 -62
rect 346 -64 348 -62
rect 361 -64 363 -62
rect 430 -64 432 -62
rect 452 -64 454 -62
rect 467 -64 469 -62
rect 536 -64 538 -62
rect 558 -64 560 -62
rect 573 -64 575 -62
rect 642 -64 644 -62
rect 664 -64 666 -62
rect 679 -64 681 -62
rect 748 -64 750 -62
rect 770 -64 772 -62
rect 785 -64 787 -62
rect 854 -64 856 -62
rect 876 -64 878 -62
rect 891 -64 893 -62
<< polyct1 >>
rect 98 1160 100 1162
rect 157 1155 159 1157
rect 167 1158 169 1160
rect 203 1155 205 1157
rect 82 1147 84 1149
rect 246 1160 248 1162
rect 213 1147 215 1149
rect 307 1155 309 1157
rect 230 1147 232 1149
rect 339 1155 341 1157
rect 367 1155 369 1157
rect 590 1154 592 1156
rect 622 1160 624 1162
rect 708 1163 710 1165
rect 317 1148 319 1150
rect 684 1155 686 1157
rect 606 1147 608 1149
rect 730 1160 732 1162
rect 719 1155 721 1157
rect 104 1079 106 1081
rect 89 1075 91 1077
rect 173 1083 175 1085
rect 125 1075 127 1077
rect 163 1075 165 1077
rect 217 1082 219 1084
rect 207 1075 209 1077
rect 229 1075 231 1077
rect 258 1076 260 1078
rect 273 1069 275 1071
rect 284 1067 286 1069
rect 323 1076 325 1078
rect 578 1075 580 1077
rect 303 1067 305 1069
rect 313 1070 315 1072
rect 630 1083 632 1085
rect 620 1075 622 1077
rect 313 1059 315 1061
rect 649 1079 651 1081
rect 739 1083 741 1085
rect 664 1075 666 1077
rect 723 1070 725 1072
rect 98 1016 100 1018
rect 157 1011 159 1013
rect 204 1017 206 1019
rect 194 1011 196 1013
rect 82 1003 84 1005
rect 172 1007 174 1009
rect 215 1019 217 1021
rect 227 1019 229 1021
rect 237 1019 239 1021
rect 265 1011 267 1013
rect 584 1019 586 1021
rect 287 1011 289 1013
rect 277 1004 279 1006
rect 520 1011 522 1013
rect 606 1016 608 1018
rect 595 1011 597 1013
rect 708 1019 710 1021
rect 642 1011 644 1013
rect 632 1003 634 1005
rect 682 1011 684 1013
rect 730 1016 732 1018
rect 719 1011 721 1013
rect 89 931 91 933
rect 173 939 175 941
rect 256 939 258 941
rect 99 928 101 930
rect 125 931 127 933
rect 163 931 165 933
rect 273 939 275 941
rect 240 926 242 928
rect 567 939 569 941
rect 283 931 285 933
rect 608 939 610 941
rect 739 939 741 941
rect 551 926 553 928
rect 598 931 600 933
rect 632 931 634 933
rect 664 931 666 933
rect 723 926 725 928
rect 87 874 89 876
rect 98 867 100 869
rect 135 867 137 869
rect 184 867 186 869
rect 145 859 147 861
rect 233 867 235 869
rect 194 859 196 861
rect 223 859 225 861
rect 273 867 275 869
rect 311 867 313 869
rect 355 867 357 869
rect 321 859 323 861
rect 377 867 379 869
rect 365 860 367 862
rect 501 867 503 869
rect 491 859 493 861
rect 540 867 542 869
rect 574 867 576 869
rect 564 859 566 861
rect 626 867 628 869
rect 656 867 658 869
rect 636 859 638 861
rect 678 867 680 869
rect 712 867 714 869
rect 668 860 670 862
rect 732 867 734 869
rect 722 859 724 861
rect 99 795 101 797
rect 89 787 91 789
rect 153 794 155 796
rect 109 787 111 789
rect 143 787 145 789
rect 185 795 187 797
rect 165 787 167 789
rect 195 787 197 789
rect 257 795 259 797
rect 247 787 249 789
rect 281 787 283 789
rect 330 795 332 797
rect 320 787 322 789
rect 456 794 458 796
rect 444 787 446 789
rect 500 795 502 797
rect 466 787 468 789
rect 510 787 512 789
rect 548 787 550 789
rect 598 795 600 797
rect 627 795 629 797
rect 588 787 590 789
rect 676 795 678 797
rect 637 787 639 789
rect 686 787 688 789
rect 723 787 725 789
rect 734 780 736 782
rect 98 728 100 730
rect 157 723 159 725
rect 189 723 191 725
rect 223 723 225 725
rect 270 728 272 730
rect 82 715 84 717
rect 213 715 215 717
rect 329 723 331 725
rect 538 723 540 725
rect 254 715 256 717
rect 581 728 583 730
rect 548 715 550 717
rect 658 723 660 725
rect 696 723 698 725
rect 722 726 724 728
rect 565 715 567 717
rect 648 715 650 717
rect 732 723 734 725
rect 102 643 104 645
rect 91 638 93 640
rect 139 643 141 645
rect 189 651 191 653
rect 179 643 181 645
rect 113 635 115 637
rect 226 643 228 645
rect 215 638 217 640
rect 544 650 546 652
rect 534 643 536 645
rect 556 643 558 645
rect 237 635 239 637
rect 584 635 586 637
rect 594 635 596 637
rect 606 635 608 637
rect 649 647 651 649
rect 739 651 741 653
rect 627 643 629 645
rect 617 637 619 639
rect 664 643 666 645
rect 723 638 725 640
rect 98 584 100 586
rect 157 579 159 581
rect 82 571 84 573
rect 172 575 174 577
rect 508 595 510 597
rect 201 579 203 581
rect 191 571 193 573
rect 508 584 510 586
rect 518 587 520 589
rect 243 579 245 581
rect 498 578 500 580
rect 537 587 539 589
rect 548 585 550 587
rect 563 578 565 580
rect 592 579 594 581
rect 614 579 616 581
rect 604 572 606 574
rect 658 579 660 581
rect 696 579 698 581
rect 648 571 650 573
rect 732 579 734 581
rect 717 575 719 577
rect 102 499 104 501
rect 91 494 93 496
rect 215 507 217 509
rect 137 499 139 501
rect 504 506 506 508
rect 113 491 115 493
rect 199 494 201 496
rect 231 500 233 502
rect 454 499 456 501
rect 482 499 484 501
rect 591 507 593 509
rect 514 499 516 501
rect 608 507 610 509
rect 575 494 577 496
rect 739 507 741 509
rect 618 499 620 501
rect 654 496 656 498
rect 664 499 666 501
rect 723 494 725 496
rect 12 332 14 334
rect 76 333 78 335
rect 86 335 88 337
rect 112 332 114 334
rect 176 333 178 335
rect 186 335 188 337
rect 212 332 214 334
rect 276 333 278 335
rect 286 335 288 337
rect 312 332 314 334
rect 376 333 378 335
rect 386 335 388 337
rect 412 332 414 334
rect 476 333 478 335
rect 486 335 488 337
rect 512 332 514 334
rect 576 333 578 335
rect 586 335 588 337
rect 612 332 614 334
rect 676 333 678 335
rect 686 335 688 337
rect 712 332 714 334
rect 776 333 778 335
rect 786 335 788 337
rect 14 249 16 251
rect 24 251 26 253
rect 88 252 90 254
rect 114 249 116 251
rect 124 251 126 253
rect 188 252 190 254
rect 214 249 216 251
rect 224 251 226 253
rect 288 252 290 254
rect 314 249 316 251
rect 324 251 326 253
rect 388 252 390 254
rect 416 249 418 251
rect 426 251 428 253
rect 490 252 492 254
rect 516 249 518 251
rect 526 251 528 253
rect 590 252 592 254
rect 616 249 618 251
rect 626 251 628 253
rect 690 252 692 254
rect 716 249 718 251
rect 726 251 728 253
rect 790 252 792 254
rect 14 191 16 193
rect 24 189 26 191
rect 88 188 90 190
rect 114 191 116 193
rect 124 190 126 192
rect 188 188 190 190
rect 214 191 216 193
rect 224 189 226 191
rect 288 188 290 190
rect 314 191 316 193
rect 324 190 326 192
rect 387 188 389 190
rect 416 191 418 193
rect 426 189 428 191
rect 490 188 492 190
rect 516 191 518 193
rect 526 190 528 192
rect 590 188 592 190
rect 616 191 618 193
rect 626 189 628 191
rect 690 188 692 190
rect 716 191 718 193
rect 726 190 728 192
rect 790 188 792 190
rect 14 105 16 107
rect 24 107 26 109
rect 88 108 90 110
rect 114 105 116 107
rect 125 107 127 109
rect 188 108 190 110
rect 214 105 216 107
rect 224 107 226 109
rect 288 108 290 110
rect 314 105 316 107
rect 324 107 326 109
rect 388 108 390 110
rect 416 105 418 107
rect 426 107 428 109
rect 490 108 492 110
rect 516 105 518 107
rect 526 107 528 109
rect 590 108 592 110
rect 616 105 618 107
rect 626 107 628 109
rect 690 108 692 110
rect 716 105 718 107
rect 726 107 728 109
rect 790 108 792 110
rect 12 44 14 46
rect 76 45 78 47
rect 86 47 88 49
rect 112 44 114 46
rect 176 45 178 47
rect 186 47 188 49
rect 212 44 214 46
rect 276 45 278 47
rect 286 47 288 49
rect 312 44 314 46
rect 376 45 378 47
rect 386 47 388 49
rect 412 44 414 46
rect 476 45 478 47
rect 486 47 488 49
rect 512 44 514 46
rect 576 45 578 47
rect 586 47 588 49
rect 612 44 614 46
rect 676 45 678 47
rect 686 47 688 49
rect 712 44 714 46
rect 776 45 778 47
rect 786 47 788 49
rect -5 -64 -3 -62
rect 59 -65 61 -63
rect 69 -67 71 -65
rect 101 -64 103 -62
rect 165 -65 167 -63
rect 175 -67 177 -65
rect 207 -64 209 -62
rect 271 -65 273 -63
rect 281 -67 283 -65
rect 313 -64 315 -62
rect 377 -65 379 -63
rect 387 -67 389 -65
rect 419 -64 421 -62
rect 483 -65 485 -63
rect 493 -67 495 -65
rect 525 -64 527 -62
rect 589 -65 591 -63
rect 599 -67 601 -65
rect 631 -64 633 -62
rect 695 -65 697 -63
rect 705 -67 707 -65
rect 737 -64 739 -62
rect 801 -65 803 -63
rect 811 -67 813 -65
rect 843 -64 845 -62
rect 907 -65 909 -63
rect 917 -67 919 -65
<< ndifct0 >>
rect 96 1172 98 1174
rect 82 1164 84 1166
rect 108 1169 110 1171
rect 172 1169 174 1171
rect 216 1171 218 1173
rect 244 1172 246 1174
rect 230 1164 232 1166
rect 256 1169 258 1171
rect 568 1171 570 1173
rect 374 1167 376 1169
rect 620 1172 622 1174
rect 590 1168 592 1170
rect 606 1164 608 1166
rect 632 1169 634 1171
rect 717 1178 719 1180
rect 717 1171 719 1173
rect 691 1167 693 1169
rect 737 1178 739 1180
rect 132 1063 134 1065
rect 104 1059 106 1061
rect 176 1059 178 1061
rect 104 1052 106 1054
rect 227 1058 229 1060
rect 258 1058 260 1060
rect 300 1058 302 1060
rect 571 1063 573 1065
rect 633 1059 635 1061
rect 649 1059 651 1061
rect 649 1052 651 1054
rect 713 1061 715 1063
rect 739 1066 741 1068
rect 725 1058 727 1060
rect 96 1028 98 1030
rect 82 1020 84 1022
rect 108 1025 110 1027
rect 172 1034 174 1036
rect 172 1027 174 1029
rect 267 1028 269 1030
rect 593 1034 595 1036
rect 593 1027 595 1029
rect 527 1023 529 1025
rect 613 1034 615 1036
rect 629 1027 631 1029
rect 717 1034 719 1036
rect 717 1027 719 1029
rect 689 1023 691 1025
rect 737 1034 739 1036
rect 104 917 106 919
rect 132 919 134 921
rect 176 915 178 917
rect 230 917 232 919
rect 256 922 258 924
rect 242 914 244 916
rect 270 915 272 917
rect 541 917 543 919
rect 567 922 569 924
rect 553 914 555 916
rect 625 922 627 924
rect 611 915 613 917
rect 636 913 638 915
rect 646 921 648 923
rect 646 914 648 916
rect 666 914 668 916
rect 713 917 715 919
rect 739 922 741 924
rect 725 914 727 916
rect 83 889 85 891
rect 148 883 150 885
rect 197 883 199 885
rect 220 883 222 885
rect 280 879 282 881
rect 324 883 326 885
rect 375 884 377 886
rect 488 883 490 885
rect 561 883 563 885
rect 547 879 549 881
rect 711 891 713 892
rect 639 883 641 885
rect 658 884 660 886
rect 163 770 165 772
rect 182 771 184 773
rect 110 764 112 765
rect 274 775 276 777
rect 260 771 262 773
rect 333 771 335 773
rect 446 770 448 772
rect 497 771 499 773
rect 541 775 543 777
rect 601 771 603 773
rect 624 771 626 773
rect 673 771 675 773
rect 738 765 740 767
rect 96 740 98 742
rect 82 732 84 734
rect 108 737 110 739
rect 155 740 157 742
rect 175 740 177 742
rect 175 733 177 735
rect 185 741 187 743
rect 210 739 212 741
rect 196 732 198 734
rect 268 740 270 742
rect 254 732 256 734
rect 280 737 282 739
rect 336 735 338 737
rect 551 739 553 741
rect 579 740 581 742
rect 565 732 567 734
rect 591 737 593 739
rect 645 739 647 741
rect 689 735 691 737
rect 717 737 719 739
rect 84 620 86 622
rect 132 631 134 633
rect 104 627 106 629
rect 104 620 106 622
rect 192 627 194 629
rect 208 620 210 622
rect 228 627 230 629
rect 228 620 230 622
rect 554 626 556 628
rect 649 627 651 629
rect 649 620 651 622
rect 713 629 715 631
rect 739 634 741 636
rect 725 626 727 628
rect 96 596 98 598
rect 82 588 84 590
rect 108 593 110 595
rect 172 602 174 604
rect 172 595 174 597
rect 188 595 190 597
rect 250 591 252 593
rect 521 596 523 598
rect 563 596 565 598
rect 594 596 596 598
rect 717 602 719 604
rect 645 595 647 597
rect 717 595 719 597
rect 689 591 691 593
rect 84 476 86 478
rect 130 487 132 489
rect 104 483 106 485
rect 104 476 106 478
rect 189 485 191 487
rect 215 490 217 492
rect 231 486 233 488
rect 201 482 203 484
rect 447 487 449 489
rect 253 483 255 485
rect 565 485 567 487
rect 591 490 593 492
rect 577 482 579 484
rect 605 483 607 485
rect 649 485 651 487
rect 713 485 715 487
rect 739 490 741 492
rect 725 482 727 484
rect 9 342 11 344
rect 20 347 22 349
rect 30 342 32 344
rect 50 347 52 349
rect 82 355 84 357
rect 60 349 62 351
rect 70 344 72 346
rect 93 344 95 346
rect 109 342 111 344
rect 120 347 122 349
rect 130 342 132 344
rect 150 347 152 349
rect 182 355 184 357
rect 160 349 162 351
rect 170 344 172 346
rect 193 344 195 346
rect 209 342 211 344
rect 220 347 222 349
rect 230 342 232 344
rect 250 347 252 349
rect 282 355 284 357
rect 260 349 262 351
rect 270 344 272 346
rect 293 344 295 346
rect 309 342 311 344
rect 320 347 322 349
rect 330 342 332 344
rect 350 347 352 349
rect 382 355 384 357
rect 360 349 362 351
rect 370 344 372 346
rect 393 344 395 346
rect 409 342 411 344
rect 420 347 422 349
rect 430 342 432 344
rect 450 347 452 349
rect 482 355 484 357
rect 460 349 462 351
rect 470 344 472 346
rect 493 344 495 346
rect 509 342 511 344
rect 520 347 522 349
rect 530 342 532 344
rect 550 347 552 349
rect 582 355 584 357
rect 560 349 562 351
rect 570 344 572 346
rect 593 344 595 346
rect 609 342 611 344
rect 620 347 622 349
rect 630 342 632 344
rect 650 347 652 349
rect 682 355 684 357
rect 660 349 662 351
rect 670 344 672 346
rect 693 344 695 346
rect 709 342 711 344
rect 720 347 722 349
rect 730 342 732 344
rect 750 347 752 349
rect 782 355 784 357
rect 760 349 762 351
rect 770 344 772 346
rect 793 344 795 346
rect 7 240 9 242
rect 30 240 32 242
rect 40 235 42 237
rect 18 229 20 231
rect 50 237 52 239
rect 70 242 72 244
rect 80 237 82 239
rect 91 242 93 244
rect 107 240 109 242
rect 130 240 132 242
rect 140 235 142 237
rect 118 229 120 231
rect 150 237 152 239
rect 170 242 172 244
rect 180 237 182 239
rect 191 242 193 244
rect 207 240 209 242
rect 230 240 232 242
rect 240 235 242 237
rect 218 229 220 231
rect 250 237 252 239
rect 270 242 272 244
rect 280 237 282 239
rect 291 242 293 244
rect 307 240 309 242
rect 330 240 332 242
rect 340 235 342 237
rect 318 229 320 231
rect 350 237 352 239
rect 370 242 372 244
rect 380 237 382 239
rect 391 242 393 244
rect 409 240 411 242
rect 432 240 434 242
rect 442 235 444 237
rect 420 229 422 231
rect 452 237 454 239
rect 472 242 474 244
rect 482 237 484 239
rect 493 242 495 244
rect 509 240 511 242
rect 532 240 534 242
rect 542 235 544 237
rect 520 229 522 231
rect 552 237 554 239
rect 572 242 574 244
rect 582 237 584 239
rect 593 242 595 244
rect 609 240 611 242
rect 632 240 634 242
rect 642 235 644 237
rect 620 229 622 231
rect 652 237 654 239
rect 672 242 674 244
rect 682 237 684 239
rect 693 242 695 244
rect 709 240 711 242
rect 732 240 734 242
rect 742 235 744 237
rect 720 229 722 231
rect 752 237 754 239
rect 772 242 774 244
rect 782 237 784 239
rect 793 242 795 244
rect 18 211 20 213
rect 7 200 9 202
rect 40 205 42 207
rect 30 200 32 202
rect 50 203 52 205
rect 70 198 72 200
rect 80 203 82 205
rect 118 211 120 213
rect 91 198 93 200
rect 107 200 109 202
rect 140 205 142 207
rect 130 200 132 202
rect 150 203 152 205
rect 170 198 172 200
rect 180 203 182 205
rect 218 211 220 213
rect 191 198 193 200
rect 207 200 209 202
rect 240 205 242 207
rect 230 200 232 202
rect 250 203 252 205
rect 270 198 272 200
rect 280 203 282 205
rect 318 211 320 213
rect 291 198 293 200
rect 307 200 309 202
rect 340 205 342 207
rect 330 200 332 202
rect 350 203 352 205
rect 370 198 372 200
rect 380 203 382 205
rect 420 211 422 213
rect 391 198 393 200
rect 409 200 411 202
rect 442 205 444 207
rect 432 200 434 202
rect 452 203 454 205
rect 472 198 474 200
rect 482 203 484 205
rect 520 211 522 213
rect 493 198 495 200
rect 509 200 511 202
rect 542 205 544 207
rect 532 200 534 202
rect 552 203 554 205
rect 572 198 574 200
rect 582 203 584 205
rect 620 211 622 213
rect 593 198 595 200
rect 609 200 611 202
rect 642 205 644 207
rect 632 200 634 202
rect 652 203 654 205
rect 672 198 674 200
rect 682 203 684 205
rect 720 211 722 213
rect 693 198 695 200
rect 709 200 711 202
rect 742 205 744 207
rect 732 200 734 202
rect 752 203 754 205
rect 772 198 774 200
rect 782 203 784 205
rect 793 198 795 200
rect 7 96 9 98
rect 30 96 32 98
rect 40 91 42 93
rect 18 85 20 87
rect 50 93 52 95
rect 70 98 72 100
rect 80 93 82 95
rect 91 98 93 100
rect 107 96 109 98
rect 130 96 132 98
rect 140 91 142 93
rect 118 85 120 87
rect 150 93 152 95
rect 170 98 172 100
rect 180 93 182 95
rect 191 98 193 100
rect 207 96 209 98
rect 230 96 232 98
rect 240 91 242 93
rect 218 85 220 87
rect 250 93 252 95
rect 270 98 272 100
rect 280 93 282 95
rect 291 98 293 100
rect 307 96 309 98
rect 330 96 332 98
rect 340 91 342 93
rect 318 85 320 87
rect 350 93 352 95
rect 370 98 372 100
rect 380 93 382 95
rect 391 98 393 100
rect 409 96 411 98
rect 432 96 434 98
rect 442 91 444 93
rect 420 85 422 87
rect 452 93 454 95
rect 472 98 474 100
rect 482 93 484 95
rect 493 98 495 100
rect 509 96 511 98
rect 532 96 534 98
rect 542 91 544 93
rect 520 85 522 87
rect 552 93 554 95
rect 572 98 574 100
rect 582 93 584 95
rect 593 98 595 100
rect 609 96 611 98
rect 632 96 634 98
rect 642 91 644 93
rect 620 85 622 87
rect 652 93 654 95
rect 672 98 674 100
rect 682 93 684 95
rect 693 98 695 100
rect 709 96 711 98
rect 732 96 734 98
rect 742 91 744 93
rect 720 85 722 87
rect 752 93 754 95
rect 772 98 774 100
rect 782 93 784 95
rect 793 98 795 100
rect 9 54 11 56
rect 20 59 22 61
rect 30 54 32 56
rect 50 59 52 61
rect 82 67 84 69
rect 60 61 62 63
rect 70 56 72 58
rect 93 56 95 58
rect 109 54 111 56
rect 120 59 122 61
rect 130 54 132 56
rect 150 59 152 61
rect 182 67 184 69
rect 160 61 162 63
rect 170 56 172 58
rect 193 56 195 58
rect 209 54 211 56
rect 220 59 222 61
rect 230 54 232 56
rect 250 59 252 61
rect 282 67 284 69
rect 260 61 262 63
rect 270 56 272 58
rect 293 56 295 58
rect 309 54 311 56
rect 320 59 322 61
rect 330 54 332 56
rect 350 59 352 61
rect 382 67 384 69
rect 360 61 362 63
rect 370 56 372 58
rect 393 56 395 58
rect 409 54 411 56
rect 420 59 422 61
rect 430 54 432 56
rect 450 59 452 61
rect 482 67 484 69
rect 460 61 462 63
rect 470 56 472 58
rect 493 56 495 58
rect 509 54 511 56
rect 520 59 522 61
rect 530 54 532 56
rect 550 59 552 61
rect 582 67 584 69
rect 560 61 562 63
rect 570 56 572 58
rect 593 56 595 58
rect 609 54 611 56
rect 620 59 622 61
rect 630 54 632 56
rect 650 59 652 61
rect 682 67 684 69
rect 660 61 662 63
rect 670 56 672 58
rect 693 56 695 58
rect 709 54 711 56
rect 720 59 722 61
rect 730 54 732 56
rect 750 59 752 61
rect 782 67 784 69
rect 760 61 762 63
rect 770 56 772 58
rect 793 56 795 58
rect -8 -74 -6 -72
rect 3 -79 5 -77
rect 13 -74 15 -72
rect 33 -79 35 -77
rect 53 -76 55 -74
rect 43 -81 45 -79
rect 76 -76 78 -74
rect 98 -74 100 -72
rect 65 -87 67 -85
rect 109 -79 111 -77
rect 119 -74 121 -72
rect 139 -79 141 -77
rect 159 -76 161 -74
rect 149 -81 151 -79
rect 182 -76 184 -74
rect 204 -74 206 -72
rect 171 -87 173 -85
rect 215 -79 217 -77
rect 225 -74 227 -72
rect 245 -79 247 -77
rect 265 -76 267 -74
rect 255 -81 257 -79
rect 288 -76 290 -74
rect 310 -74 312 -72
rect 277 -87 279 -85
rect 321 -79 323 -77
rect 331 -74 333 -72
rect 351 -79 353 -77
rect 371 -76 373 -74
rect 361 -81 363 -79
rect 394 -76 396 -74
rect 416 -74 418 -72
rect 383 -87 385 -85
rect 427 -79 429 -77
rect 437 -74 439 -72
rect 457 -79 459 -77
rect 477 -76 479 -74
rect 467 -81 469 -79
rect 500 -76 502 -74
rect 522 -74 524 -72
rect 489 -87 491 -85
rect 533 -79 535 -77
rect 543 -74 545 -72
rect 563 -79 565 -77
rect 583 -76 585 -74
rect 573 -81 575 -79
rect 606 -76 608 -74
rect 628 -74 630 -72
rect 595 -87 597 -85
rect 639 -79 641 -77
rect 649 -74 651 -72
rect 669 -79 671 -77
rect 689 -76 691 -74
rect 679 -81 681 -79
rect 712 -76 714 -74
rect 734 -74 736 -72
rect 701 -87 703 -85
rect 745 -79 747 -77
rect 755 -74 757 -72
rect 775 -79 777 -77
rect 795 -76 797 -74
rect 785 -81 787 -79
rect 818 -76 820 -74
rect 840 -74 842 -72
rect 807 -87 809 -85
rect 851 -79 853 -77
rect 861 -74 863 -72
rect 881 -79 883 -77
rect 901 -76 903 -74
rect 891 -81 893 -79
rect 924 -76 926 -74
rect 913 -87 915 -85
<< ndifct1 >>
rect 136 1181 138 1183
rect 118 1171 120 1173
rect 150 1181 152 1183
rect 197 1181 199 1183
rect 161 1172 163 1174
rect 284 1181 286 1183
rect 186 1169 188 1171
rect 266 1171 268 1173
rect 306 1172 308 1174
rect 338 1181 340 1183
rect 660 1181 662 1183
rect 360 1164 362 1166
rect 579 1164 581 1166
rect 642 1171 644 1173
rect 677 1164 679 1166
rect 727 1171 729 1173
rect 85 1058 87 1060
rect 118 1066 120 1068
rect 146 1061 148 1063
rect 190 1065 192 1067
rect 268 1058 270 1060
rect 290 1058 292 1060
rect 157 1049 159 1051
rect 585 1066 587 1068
rect 603 1061 605 1063
rect 201 1049 203 1051
rect 279 1049 281 1051
rect 614 1049 616 1051
rect 668 1058 670 1060
rect 703 1059 705 1061
rect 685 1049 687 1051
rect 136 1037 138 1039
rect 118 1027 120 1029
rect 153 1028 155 1030
rect 211 1037 213 1039
rect 233 1037 235 1039
rect 293 1037 295 1039
rect 222 1028 224 1030
rect 244 1028 246 1030
rect 304 1021 306 1023
rect 513 1020 515 1022
rect 603 1027 605 1029
rect 648 1037 650 1039
rect 659 1025 661 1027
rect 675 1020 677 1022
rect 727 1027 729 1029
rect 93 914 95 916
rect 118 922 120 924
rect 146 917 148 919
rect 82 905 84 907
rect 220 915 222 917
rect 300 917 302 919
rect 157 905 159 907
rect 202 905 204 907
rect 531 915 533 917
rect 581 917 583 919
rect 289 905 291 907
rect 513 905 515 907
rect 592 905 594 907
rect 656 922 658 924
rect 703 915 705 917
rect 685 905 687 907
rect 129 893 131 895
rect 178 893 180 895
rect 105 883 107 885
rect 118 881 120 883
rect 239 893 241 895
rect 305 893 307 895
rect 167 881 169 883
rect 349 893 351 895
rect 507 893 509 895
rect 250 881 252 883
rect 266 876 268 878
rect 294 881 296 883
rect 338 877 340 879
rect 580 893 582 895
rect 620 893 622 895
rect 684 893 686 895
rect 518 881 520 883
rect 533 876 535 878
rect 711 892 713 893
rect 591 881 593 883
rect 609 881 611 883
rect 695 877 697 879
rect 736 884 738 886
rect 85 770 87 772
rect 126 777 128 779
rect 212 773 214 775
rect 230 773 232 775
rect 110 763 112 764
rect 288 778 290 780
rect 303 773 305 775
rect 137 761 139 763
rect 201 761 203 763
rect 241 761 243 763
rect 483 777 485 779
rect 527 773 529 775
rect 555 778 557 780
rect 571 773 573 775
rect 314 761 316 763
rect 472 761 474 763
rect 654 773 656 775
rect 516 761 518 763
rect 582 761 584 763
rect 703 773 705 775
rect 716 771 718 773
rect 643 761 645 763
rect 692 761 694 763
rect 136 749 138 751
rect 118 739 120 741
rect 165 732 167 734
rect 229 749 231 751
rect 308 749 310 751
rect 532 749 534 751
rect 240 737 242 739
rect 290 739 292 741
rect 619 749 621 751
rect 664 749 666 751
rect 322 732 324 734
rect 521 737 523 739
rect 601 739 603 741
rect 739 749 741 751
rect 675 737 677 739
rect 703 732 705 734
rect 728 740 730 742
rect 94 627 96 629
rect 146 634 148 636
rect 162 629 164 631
rect 517 633 519 635
rect 173 617 175 619
rect 218 627 220 629
rect 577 626 579 628
rect 599 626 601 628
rect 528 617 530 619
rect 588 617 590 619
rect 610 617 612 619
rect 668 626 670 628
rect 703 627 705 629
rect 685 617 687 619
rect 136 605 138 607
rect 118 595 120 597
rect 153 596 155 598
rect 207 605 209 607
rect 542 605 544 607
rect 620 605 622 607
rect 218 593 220 595
rect 236 588 238 590
rect 664 605 666 607
rect 531 596 533 598
rect 553 596 555 598
rect 631 589 633 591
rect 675 593 677 595
rect 703 588 705 590
rect 736 596 738 598
rect 94 483 96 485
rect 144 490 146 492
rect 179 483 181 485
rect 242 490 244 492
rect 461 490 463 492
rect 161 473 163 475
rect 483 473 485 475
rect 515 482 517 484
rect 555 483 557 485
rect 635 485 637 487
rect 537 473 539 475
rect 660 482 662 484
rect 624 473 626 475
rect 671 473 673 475
rect 703 483 705 485
rect 685 473 687 475
rect 40 347 42 349
rect 140 347 142 349
rect 240 347 242 349
rect 340 347 342 349
rect 440 347 442 349
rect 540 347 542 349
rect 640 347 642 349
rect 740 347 742 349
rect 60 237 62 239
rect 160 237 162 239
rect 260 237 262 239
rect 360 237 362 239
rect 462 237 464 239
rect 562 237 564 239
rect 662 237 664 239
rect 762 237 764 239
rect 60 203 62 205
rect 160 203 162 205
rect 260 203 262 205
rect 360 203 362 205
rect 462 203 464 205
rect 562 203 564 205
rect 662 203 664 205
rect 762 203 764 205
rect 60 93 62 95
rect 160 93 162 95
rect 260 93 262 95
rect 360 93 362 95
rect 462 93 464 95
rect 562 93 564 95
rect 662 93 664 95
rect 762 93 764 95
rect 40 59 42 61
rect 140 59 142 61
rect 240 59 242 61
rect 340 59 342 61
rect 440 59 442 61
rect 540 59 542 61
rect 640 59 642 61
rect 740 59 742 61
rect 23 -79 25 -77
rect 129 -79 131 -77
rect 235 -79 237 -77
rect 341 -79 343 -77
rect 447 -79 449 -77
rect 553 -79 555 -77
rect 659 -79 661 -77
rect 765 -79 767 -77
rect 871 -79 873 -77
<< ntiect1 >>
rect 116 1121 118 1123
rect 187 1121 189 1123
rect 264 1121 266 1123
rect 361 1121 363 1123
rect 373 1121 375 1123
rect 588 1121 590 1123
rect 640 1121 642 1123
rect 678 1121 680 1123
rect 690 1121 692 1123
rect 119 1109 121 1111
rect 131 1109 133 1111
rect 147 1109 149 1111
rect 235 1109 237 1111
rect 301 1109 303 1111
rect 323 1109 325 1111
rect 572 1109 574 1111
rect 584 1109 586 1111
rect 604 1109 606 1111
rect 705 1109 707 1111
rect 116 977 118 979
rect 259 977 261 979
rect 514 977 516 979
rect 526 977 528 979
rect 658 977 660 979
rect 676 977 678 979
rect 688 977 690 979
rect 119 965 121 967
rect 131 965 133 967
rect 147 965 149 967
rect 222 965 224 967
rect 299 965 301 967
rect 533 965 535 967
rect 582 965 584 967
rect 626 965 628 967
rect 634 965 636 967
rect 705 965 707 967
rect 84 833 86 835
rect 92 833 94 835
rect 119 833 121 835
rect 168 833 170 835
rect 249 833 251 835
rect 267 833 269 835
rect 279 833 281 835
rect 295 833 297 835
rect 383 833 385 835
rect 517 833 519 835
rect 534 833 536 835
rect 546 833 548 835
rect 590 833 592 835
rect 610 833 612 835
rect 650 833 652 835
rect 171 821 173 823
rect 211 821 213 823
rect 231 821 233 823
rect 275 821 277 823
rect 287 821 289 823
rect 304 821 306 823
rect 438 821 440 823
rect 526 821 528 823
rect 542 821 544 823
rect 554 821 556 823
rect 572 821 574 823
rect 653 821 655 823
rect 702 821 704 823
rect 729 821 731 823
rect 737 821 739 823
rect 116 689 118 691
rect 187 689 189 691
rect 195 689 197 691
rect 239 689 241 691
rect 288 689 290 691
rect 323 689 325 691
rect 335 689 337 691
rect 522 689 524 691
rect 599 689 601 691
rect 674 689 676 691
rect 690 689 692 691
rect 702 689 704 691
rect 133 677 135 679
rect 145 677 147 679
rect 163 677 165 679
rect 562 677 564 679
rect 705 677 707 679
rect 116 545 118 547
rect 217 545 219 547
rect 237 545 239 547
rect 249 545 251 547
rect 498 545 500 547
rect 520 545 522 547
rect 586 545 588 547
rect 674 545 676 547
rect 690 545 692 547
rect 702 545 704 547
rect 131 533 133 535
rect 143 533 145 535
rect 181 533 183 535
rect 233 533 235 535
rect 448 533 450 535
rect 460 533 462 535
rect 557 533 559 535
rect 634 533 636 535
rect 705 533 707 535
rect 8 298 10 300
rect 108 298 110 300
rect 208 298 210 300
rect 308 298 310 300
rect 408 298 410 300
rect 508 298 510 300
rect 608 298 610 300
rect 708 298 710 300
rect 92 286 94 288
rect 192 286 194 288
rect 292 286 294 288
rect 392 286 394 288
rect 494 286 496 288
rect 594 286 596 288
rect 694 286 696 288
rect 794 286 796 288
rect 92 154 94 156
rect 192 154 194 156
rect 292 154 294 156
rect 392 154 394 156
rect 494 154 496 156
rect 594 154 596 156
rect 694 154 696 156
rect 794 154 796 156
rect 92 142 94 144
rect 192 142 194 144
rect 292 142 294 144
rect 392 142 394 144
rect 494 142 496 144
rect 594 142 596 144
rect 694 142 696 144
rect 794 142 796 144
rect 8 10 10 12
rect 108 10 110 12
rect 208 10 210 12
rect 308 10 310 12
rect 408 10 410 12
rect 508 10 510 12
rect 608 10 610 12
rect 708 10 710 12
rect -9 -30 -7 -28
rect 97 -30 99 -28
rect 203 -30 205 -28
rect 309 -30 311 -28
rect 415 -30 417 -28
rect 521 -30 523 -28
rect 627 -30 629 -28
rect 733 -30 735 -28
rect 839 -30 841 -28
<< ptiect1 >>
rect 83 1181 85 1183
rect 171 1181 173 1183
rect 187 1181 189 1183
rect 231 1181 233 1183
rect 361 1181 363 1183
rect 373 1181 375 1183
rect 569 1181 571 1183
rect 589 1181 591 1183
rect 607 1181 609 1183
rect 678 1181 680 1183
rect 690 1181 692 1183
rect 702 1181 704 1183
rect 119 1049 121 1051
rect 131 1049 133 1051
rect 147 1049 149 1051
rect 191 1049 193 1051
rect 323 1049 325 1051
rect 572 1049 574 1051
rect 584 1049 586 1051
rect 604 1049 606 1051
rect 738 1049 740 1051
rect 83 1037 85 1039
rect 195 1037 197 1039
rect 303 1037 305 1039
rect 514 1037 516 1039
rect 526 1037 528 1039
rect 578 1037 580 1039
rect 658 1037 660 1039
rect 676 1037 678 1039
rect 688 1037 690 1039
rect 702 1037 704 1039
rect 103 905 105 907
rect 119 905 121 907
rect 131 905 133 907
rect 147 905 149 907
rect 255 905 257 907
rect 299 905 301 907
rect 566 905 568 907
rect 582 905 584 907
rect 626 905 628 907
rect 738 905 740 907
rect 119 893 121 895
rect 168 893 170 895
rect 249 893 251 895
rect 267 893 269 895
rect 279 893 281 895
rect 295 893 297 895
rect 339 893 341 895
rect 517 893 519 895
rect 534 893 536 895
rect 546 893 548 895
rect 590 893 592 895
rect 610 893 612 895
rect 694 893 696 895
rect 127 761 129 763
rect 211 761 213 763
rect 231 761 233 763
rect 275 761 277 763
rect 287 761 289 763
rect 304 761 306 763
rect 482 761 484 763
rect 526 761 528 763
rect 542 761 544 763
rect 554 761 556 763
rect 572 761 574 763
rect 653 761 655 763
rect 702 761 704 763
rect 83 749 85 751
rect 195 749 197 751
rect 239 749 241 751
rect 255 749 257 751
rect 323 749 325 751
rect 335 749 337 751
rect 522 749 524 751
rect 566 749 568 751
rect 674 749 676 751
rect 690 749 692 751
rect 702 749 704 751
rect 718 749 720 751
rect 119 617 121 619
rect 133 617 135 619
rect 145 617 147 619
rect 163 617 165 619
rect 243 617 245 619
rect 518 617 520 619
rect 626 617 628 619
rect 738 617 740 619
rect 83 605 85 607
rect 217 605 219 607
rect 237 605 239 607
rect 249 605 251 607
rect 498 605 500 607
rect 630 605 632 607
rect 674 605 676 607
rect 690 605 692 607
rect 702 605 704 607
rect 119 473 121 475
rect 131 473 133 475
rect 143 473 145 475
rect 214 473 216 475
rect 232 473 234 475
rect 252 473 254 475
rect 448 473 450 475
rect 460 473 462 475
rect 590 473 592 475
rect 634 473 636 475
rect 650 473 652 475
rect 738 473 740 475
rect 8 358 10 360
rect 15 358 17 360
rect 108 358 110 360
rect 115 358 117 360
rect 208 358 210 360
rect 215 358 217 360
rect 308 358 310 360
rect 315 358 317 360
rect 408 358 410 360
rect 415 358 417 360
rect 508 358 510 360
rect 515 358 517 360
rect 608 358 610 360
rect 615 358 617 360
rect 708 358 710 360
rect 715 358 717 360
rect 85 226 87 228
rect 92 226 94 228
rect 185 226 187 228
rect 192 226 194 228
rect 285 226 287 228
rect 292 226 294 228
rect 385 226 387 228
rect 392 226 394 228
rect 487 226 489 228
rect 494 226 496 228
rect 587 226 589 228
rect 594 226 596 228
rect 687 226 689 228
rect 694 226 696 228
rect 787 226 789 228
rect 794 226 796 228
rect 85 214 87 216
rect 92 214 94 216
rect 185 214 187 216
rect 192 214 194 216
rect 285 214 287 216
rect 292 214 294 216
rect 385 214 387 216
rect 392 214 394 216
rect 487 214 489 216
rect 494 214 496 216
rect 587 214 589 216
rect 594 214 596 216
rect 687 214 689 216
rect 694 214 696 216
rect 787 214 789 216
rect 794 214 796 216
rect 85 82 87 84
rect 92 82 94 84
rect 185 82 187 84
rect 192 82 194 84
rect 285 82 287 84
rect 292 82 294 84
rect 385 82 387 84
rect 392 82 394 84
rect 487 82 489 84
rect 494 82 496 84
rect 587 82 589 84
rect 594 82 596 84
rect 687 82 689 84
rect 694 82 696 84
rect 787 82 789 84
rect 794 82 796 84
rect 8 70 10 72
rect 15 70 17 72
rect 108 70 110 72
rect 115 70 117 72
rect 208 70 210 72
rect 215 70 217 72
rect 308 70 310 72
rect 315 70 317 72
rect 408 70 410 72
rect 415 70 417 72
rect 508 70 510 72
rect 515 70 517 72
rect 608 70 610 72
rect 615 70 617 72
rect 708 70 710 72
rect 715 70 717 72
rect -9 -90 -7 -88
rect -2 -90 0 -88
rect 97 -90 99 -88
rect 104 -90 106 -88
rect 203 -90 205 -88
rect 210 -90 212 -88
rect 309 -90 311 -88
rect 316 -90 318 -88
rect 415 -90 417 -88
rect 422 -90 424 -88
rect 521 -90 523 -88
rect 528 -90 530 -88
rect 627 -90 629 -88
rect 634 -90 636 -88
rect 733 -90 735 -88
rect 740 -90 742 -88
rect 839 -90 841 -88
rect 846 -90 848 -88
<< pdifct0 >>
rect 90 1145 92 1147
rect 100 1131 102 1133
rect 116 1145 118 1147
rect 116 1138 118 1140
rect 100 1124 102 1126
rect 136 1130 138 1132
rect 172 1131 174 1133
rect 238 1145 240 1147
rect 196 1133 198 1135
rect 206 1138 208 1140
rect 206 1131 208 1133
rect 216 1131 218 1133
rect 172 1124 174 1126
rect 248 1131 250 1133
rect 264 1145 266 1147
rect 264 1138 266 1140
rect 248 1124 250 1126
rect 284 1130 286 1132
rect 300 1128 302 1130
rect 310 1131 312 1133
rect 320 1128 322 1130
rect 371 1131 373 1133
rect 569 1132 571 1134
rect 569 1125 571 1127
rect 614 1145 616 1147
rect 589 1140 591 1142
rect 589 1133 591 1135
rect 624 1131 626 1133
rect 640 1145 642 1147
rect 640 1138 642 1140
rect 624 1124 626 1126
rect 660 1130 662 1132
rect 688 1131 690 1133
rect 705 1131 707 1133
rect 705 1124 707 1126
rect 739 1131 741 1133
rect 739 1124 741 1126
rect 82 1106 84 1108
rect 82 1099 84 1101
rect 92 1099 94 1101
rect 92 1092 94 1094
rect 102 1106 104 1108
rect 102 1099 104 1101
rect 129 1099 131 1101
rect 156 1097 158 1099
rect 166 1099 168 1101
rect 166 1092 168 1094
rect 176 1099 178 1101
rect 200 1098 202 1100
rect 210 1098 212 1100
rect 210 1091 212 1093
rect 232 1097 234 1099
rect 232 1090 234 1092
rect 324 1097 326 1099
rect 324 1090 326 1092
rect 574 1099 576 1101
rect 651 1106 653 1108
rect 613 1097 615 1099
rect 623 1099 625 1101
rect 623 1092 625 1094
rect 633 1099 635 1101
rect 651 1099 653 1101
rect 661 1099 663 1101
rect 661 1092 663 1094
rect 671 1106 673 1108
rect 671 1099 673 1101
rect 685 1100 687 1102
rect 721 1106 723 1108
rect 705 1092 707 1094
rect 705 1085 707 1087
rect 721 1099 723 1101
rect 731 1085 733 1087
rect 90 1001 92 1003
rect 100 987 102 989
rect 116 1001 118 1003
rect 116 994 118 996
rect 100 980 102 982
rect 136 986 138 988
rect 150 987 152 989
rect 150 980 152 982
rect 160 994 162 996
rect 160 987 162 989
rect 170 987 172 989
rect 170 980 172 982
rect 194 987 196 989
rect 194 980 196 982
rect 218 987 220 989
rect 242 987 244 989
rect 262 996 264 998
rect 262 989 264 991
rect 284 995 286 997
rect 284 988 286 990
rect 294 988 296 990
rect 242 980 244 982
rect 524 987 526 989
rect 581 987 583 989
rect 581 980 583 982
rect 615 987 617 989
rect 629 987 631 989
rect 639 994 641 996
rect 639 987 641 989
rect 649 989 651 991
rect 615 980 617 982
rect 686 987 688 989
rect 705 987 707 989
rect 705 980 707 982
rect 739 987 741 989
rect 739 980 741 982
rect 104 962 106 964
rect 104 955 106 957
rect 129 955 131 957
rect 156 953 158 955
rect 166 955 168 957
rect 166 948 168 950
rect 176 955 178 957
rect 202 956 204 958
rect 238 962 240 964
rect 222 948 224 950
rect 222 941 224 943
rect 238 955 240 957
rect 270 955 272 957
rect 280 955 282 957
rect 280 948 282 950
rect 290 953 292 955
rect 248 941 250 943
rect 513 956 515 958
rect 549 962 551 964
rect 533 948 535 950
rect 533 941 535 943
rect 549 955 551 957
rect 559 941 561 943
rect 591 953 593 955
rect 601 955 603 957
rect 601 948 603 950
rect 611 955 613 957
rect 626 953 628 955
rect 646 953 648 955
rect 646 946 648 948
rect 666 953 668 955
rect 685 956 687 958
rect 666 946 668 948
rect 721 962 723 964
rect 705 948 707 950
rect 705 941 707 943
rect 721 955 723 957
rect 731 941 733 943
rect 83 852 85 854
rect 83 845 85 847
rect 94 852 96 854
rect 94 845 96 847
rect 105 843 107 845
rect 128 845 130 847
rect 138 850 140 852
rect 138 843 140 845
rect 148 843 150 845
rect 177 845 179 847
rect 187 850 189 852
rect 187 843 189 845
rect 197 843 199 845
rect 220 843 222 845
rect 230 850 232 852
rect 230 843 232 845
rect 240 845 242 847
rect 277 843 279 845
rect 304 845 306 847
rect 314 850 316 852
rect 314 843 316 845
rect 324 843 326 845
rect 348 844 350 846
rect 358 851 360 853
rect 358 844 360 846
rect 380 852 382 854
rect 380 845 382 847
rect 488 843 490 845
rect 498 850 500 852
rect 498 843 500 845
rect 508 845 510 847
rect 544 843 546 845
rect 561 843 563 845
rect 571 850 573 852
rect 571 843 573 845
rect 581 845 583 847
rect 619 845 621 847
rect 629 850 631 852
rect 629 843 631 845
rect 639 843 641 845
rect 653 852 655 854
rect 653 845 655 847
rect 675 851 677 853
rect 675 844 677 846
rect 685 844 687 846
rect 709 843 711 845
rect 709 836 711 838
rect 729 843 731 845
rect 729 836 731 838
rect 92 818 94 820
rect 92 811 94 813
rect 112 818 114 820
rect 112 811 114 813
rect 136 810 138 812
rect 146 810 148 812
rect 146 803 148 805
rect 168 809 170 811
rect 168 802 170 804
rect 182 811 184 813
rect 192 811 194 813
rect 192 804 194 806
rect 202 809 204 811
rect 240 809 242 811
rect 250 811 252 813
rect 250 804 252 806
rect 260 811 262 813
rect 277 811 279 813
rect 313 809 315 811
rect 323 811 325 813
rect 323 804 325 806
rect 333 811 335 813
rect 441 809 443 811
rect 441 802 443 804
rect 463 810 465 812
rect 463 803 465 805
rect 473 810 475 812
rect 497 811 499 813
rect 507 811 509 813
rect 507 804 509 806
rect 517 809 519 811
rect 544 811 546 813
rect 581 809 583 811
rect 591 811 593 813
rect 591 804 593 806
rect 601 811 603 813
rect 624 811 626 813
rect 634 811 636 813
rect 634 804 636 806
rect 644 809 646 811
rect 673 811 675 813
rect 683 811 685 813
rect 683 804 685 806
rect 693 809 695 811
rect 716 811 718 813
rect 727 809 729 811
rect 727 802 729 804
rect 738 809 740 811
rect 738 802 740 804
rect 90 713 92 715
rect 100 699 102 701
rect 116 713 118 715
rect 116 706 118 708
rect 100 692 102 694
rect 155 708 157 710
rect 136 698 138 700
rect 155 701 157 703
rect 175 708 177 710
rect 175 701 177 703
rect 195 701 197 703
rect 210 699 212 701
rect 220 706 222 708
rect 220 699 222 701
rect 230 701 232 703
rect 262 713 264 715
rect 272 699 274 701
rect 288 713 290 715
rect 288 706 290 708
rect 272 692 274 694
rect 308 698 310 700
rect 333 699 335 701
rect 573 713 575 715
rect 531 701 533 703
rect 541 706 543 708
rect 541 699 543 701
rect 551 699 553 701
rect 583 699 585 701
rect 599 713 601 715
rect 599 706 601 708
rect 583 692 585 694
rect 619 698 621 700
rect 645 699 647 701
rect 655 706 657 708
rect 655 699 657 701
rect 665 701 667 703
rect 692 699 694 701
rect 717 699 719 701
rect 717 692 719 694
rect 82 674 84 676
rect 82 667 84 669
rect 116 674 118 676
rect 116 667 118 669
rect 135 667 137 669
rect 206 674 208 676
rect 172 665 174 667
rect 182 667 184 669
rect 182 660 184 662
rect 192 667 194 669
rect 206 667 208 669
rect 240 674 242 676
rect 579 674 581 676
rect 240 667 242 669
rect 527 666 529 668
rect 537 666 539 668
rect 537 659 539 661
rect 559 665 561 667
rect 559 658 561 660
rect 579 667 581 669
rect 603 667 605 669
rect 627 674 629 676
rect 627 667 629 669
rect 651 674 653 676
rect 651 667 653 669
rect 661 667 663 669
rect 661 660 663 662
rect 671 674 673 676
rect 671 667 673 669
rect 685 668 687 670
rect 721 674 723 676
rect 705 660 707 662
rect 705 653 707 655
rect 721 667 723 669
rect 731 653 733 655
rect 90 569 92 571
rect 100 555 102 557
rect 116 569 118 571
rect 116 562 118 564
rect 100 548 102 550
rect 136 554 138 556
rect 150 555 152 557
rect 150 548 152 550
rect 160 562 162 564
rect 160 555 162 557
rect 170 555 172 557
rect 188 555 190 557
rect 198 562 200 564
rect 198 555 200 557
rect 208 557 210 559
rect 170 548 172 550
rect 247 555 249 557
rect 497 564 499 566
rect 497 557 499 559
rect 589 564 591 566
rect 589 557 591 559
rect 611 563 613 565
rect 611 556 613 558
rect 621 556 623 558
rect 645 555 647 557
rect 655 562 657 564
rect 655 555 657 557
rect 665 557 667 559
rect 692 555 694 557
rect 719 555 721 557
rect 719 548 721 550
rect 729 562 731 564
rect 729 555 731 557
rect 739 555 741 557
rect 739 548 741 550
rect 82 530 84 532
rect 82 523 84 525
rect 116 530 118 532
rect 116 523 118 525
rect 133 523 135 525
rect 161 524 163 526
rect 197 530 199 532
rect 181 516 183 518
rect 181 509 183 511
rect 197 523 199 525
rect 232 521 234 523
rect 232 514 234 516
rect 207 509 209 511
rect 252 529 254 531
rect 252 522 254 524
rect 450 523 452 525
rect 501 526 503 528
rect 511 523 513 525
rect 521 526 523 528
rect 537 524 539 526
rect 573 530 575 532
rect 557 516 559 518
rect 557 509 559 511
rect 573 523 575 525
rect 649 530 651 532
rect 605 523 607 525
rect 615 523 617 525
rect 615 516 617 518
rect 625 521 627 523
rect 583 509 585 511
rect 649 523 651 525
rect 685 524 687 526
rect 721 530 723 532
rect 705 516 707 518
rect 705 509 707 511
rect 721 523 723 525
rect 731 509 733 511
rect 7 316 9 318
rect 18 308 20 310
rect 28 316 30 318
rect 52 323 54 325
rect 70 323 72 325
rect 93 315 95 317
rect 62 307 64 309
rect 81 307 83 309
rect 118 308 120 310
rect 128 316 130 318
rect 152 323 154 325
rect 170 323 172 325
rect 193 315 195 317
rect 207 316 209 318
rect 162 307 164 309
rect 181 307 183 309
rect 218 308 220 310
rect 228 316 230 318
rect 252 323 254 325
rect 270 323 272 325
rect 293 315 295 317
rect 307 316 309 318
rect 262 307 264 309
rect 281 307 283 309
rect 318 308 320 310
rect 328 316 330 318
rect 352 323 354 325
rect 370 323 372 325
rect 393 315 395 317
rect 407 316 409 318
rect 362 307 364 309
rect 381 307 383 309
rect 418 308 420 310
rect 428 316 430 318
rect 452 323 454 325
rect 470 323 472 325
rect 493 315 495 317
rect 507 316 509 318
rect 462 307 464 309
rect 481 307 483 309
rect 518 308 520 310
rect 528 316 530 318
rect 552 323 554 325
rect 570 323 572 325
rect 593 315 595 317
rect 607 316 609 318
rect 562 307 564 309
rect 581 307 583 309
rect 618 308 620 310
rect 628 316 630 318
rect 652 323 654 325
rect 670 323 672 325
rect 693 315 695 317
rect 707 316 709 318
rect 662 307 664 309
rect 681 307 683 309
rect 718 308 720 310
rect 728 316 730 318
rect 752 323 754 325
rect 770 323 772 325
rect 793 315 795 317
rect 762 307 764 309
rect 781 307 783 309
rect 19 277 21 279
rect 38 277 40 279
rect 7 269 9 271
rect 30 261 32 263
rect 48 261 50 263
rect 72 268 74 270
rect 82 276 84 278
rect 119 277 121 279
rect 138 277 140 279
rect 93 268 95 270
rect 107 269 109 271
rect 130 261 132 263
rect 148 261 150 263
rect 172 268 174 270
rect 182 276 184 278
rect 219 277 221 279
rect 238 277 240 279
rect 193 268 195 270
rect 207 269 209 271
rect 230 261 232 263
rect 248 261 250 263
rect 272 268 274 270
rect 282 276 284 278
rect 319 277 321 279
rect 338 277 340 279
rect 293 269 295 271
rect 307 269 309 271
rect 330 261 332 263
rect 348 261 350 263
rect 372 268 374 270
rect 382 276 384 278
rect 421 277 423 279
rect 440 277 442 279
rect 393 268 395 270
rect 409 269 411 271
rect 432 261 434 263
rect 450 261 452 263
rect 474 268 476 270
rect 484 276 486 278
rect 521 277 523 279
rect 540 277 542 279
rect 495 269 497 271
rect 509 269 511 271
rect 532 261 534 263
rect 550 261 552 263
rect 574 268 576 270
rect 584 276 586 278
rect 621 277 623 279
rect 640 277 642 279
rect 595 268 597 270
rect 609 269 611 271
rect 632 261 634 263
rect 650 261 652 263
rect 674 268 676 270
rect 684 276 686 278
rect 721 277 723 279
rect 740 277 742 279
rect 695 269 697 271
rect 709 269 711 271
rect 732 261 734 263
rect 750 261 752 263
rect 774 268 776 270
rect 784 276 786 278
rect 795 268 797 270
rect 7 171 9 173
rect 30 179 32 181
rect 19 163 21 165
rect 38 163 40 165
rect 48 179 50 181
rect 72 172 74 174
rect 93 172 95 174
rect 107 171 109 173
rect 82 164 84 166
rect 130 179 132 181
rect 119 163 121 165
rect 138 163 140 165
rect 148 179 150 181
rect 172 172 174 174
rect 193 172 195 174
rect 207 171 209 173
rect 182 164 184 166
rect 230 179 232 181
rect 219 163 221 165
rect 238 163 240 165
rect 248 179 250 181
rect 272 172 274 174
rect 293 172 295 174
rect 307 171 309 173
rect 282 164 284 166
rect 330 179 332 181
rect 319 163 321 165
rect 338 163 340 165
rect 348 179 350 181
rect 372 172 374 174
rect 393 172 395 174
rect 409 171 411 173
rect 382 164 384 166
rect 432 179 434 181
rect 421 163 423 165
rect 440 163 442 165
rect 450 179 452 181
rect 474 172 476 174
rect 495 172 497 174
rect 509 171 511 173
rect 484 164 486 166
rect 532 179 534 181
rect 521 163 523 165
rect 540 163 542 165
rect 550 179 552 181
rect 574 172 576 174
rect 595 172 597 174
rect 609 171 611 173
rect 584 164 586 166
rect 632 179 634 181
rect 621 163 623 165
rect 640 163 642 165
rect 650 179 652 181
rect 674 172 676 174
rect 695 172 697 174
rect 709 171 711 173
rect 684 164 686 166
rect 732 179 734 181
rect 721 163 723 165
rect 740 163 742 165
rect 750 179 752 181
rect 774 172 776 174
rect 795 172 797 174
rect 784 164 786 166
rect 19 133 21 135
rect 38 133 40 135
rect 7 125 9 127
rect 30 117 32 119
rect 48 117 50 119
rect 72 124 74 126
rect 82 132 84 134
rect 119 133 121 135
rect 138 133 140 135
rect 93 124 95 126
rect 107 125 109 127
rect 130 117 132 119
rect 148 117 150 119
rect 172 124 174 126
rect 182 132 184 134
rect 219 133 221 135
rect 238 133 240 135
rect 193 124 195 126
rect 207 125 209 127
rect 230 117 232 119
rect 248 117 250 119
rect 272 124 274 126
rect 282 132 284 134
rect 319 133 321 135
rect 338 133 340 135
rect 293 124 295 126
rect 307 125 309 127
rect 330 117 332 119
rect 348 117 350 119
rect 372 124 374 126
rect 382 132 384 134
rect 421 133 423 135
rect 440 133 442 135
rect 393 124 395 126
rect 409 125 411 127
rect 432 117 434 119
rect 450 117 452 119
rect 474 124 476 126
rect 484 132 486 134
rect 521 133 523 135
rect 540 133 542 135
rect 495 124 497 126
rect 509 125 511 127
rect 532 117 534 119
rect 550 117 552 119
rect 574 124 576 126
rect 584 132 586 134
rect 621 133 623 135
rect 640 133 642 135
rect 595 124 597 126
rect 609 125 611 127
rect 632 117 634 119
rect 650 117 652 119
rect 674 124 676 126
rect 684 132 686 134
rect 721 133 723 135
rect 740 133 742 135
rect 695 124 697 126
rect 709 125 711 127
rect 732 117 734 119
rect 750 117 752 119
rect 774 124 776 126
rect 784 132 786 134
rect 795 124 797 126
rect 7 28 9 30
rect 18 20 20 22
rect 28 28 30 30
rect 52 35 54 37
rect 70 35 72 37
rect 93 27 95 29
rect 62 19 64 21
rect 81 19 83 21
rect 118 20 120 22
rect 128 28 130 30
rect 152 35 154 37
rect 170 35 172 37
rect 193 27 195 29
rect 207 28 209 30
rect 162 19 164 21
rect 181 19 183 21
rect 218 20 220 22
rect 228 28 230 30
rect 252 35 254 37
rect 270 35 272 37
rect 293 27 295 29
rect 307 28 309 30
rect 262 19 264 21
rect 281 19 283 21
rect 318 20 320 22
rect 328 28 330 30
rect 352 35 354 37
rect 370 35 372 37
rect 393 27 395 29
rect 407 28 409 30
rect 362 19 364 21
rect 381 19 383 21
rect 418 20 420 22
rect 428 28 430 30
rect 452 35 454 37
rect 470 35 472 37
rect 493 27 495 29
rect 507 28 509 30
rect 462 19 464 21
rect 481 19 483 21
rect 518 20 520 22
rect 528 28 530 30
rect 552 35 554 37
rect 570 35 572 37
rect 593 27 595 29
rect 607 28 609 30
rect 562 19 564 21
rect 581 19 583 21
rect 618 20 620 22
rect 628 28 630 30
rect 652 35 654 37
rect 670 35 672 37
rect 693 27 695 29
rect 707 28 709 30
rect 662 19 664 21
rect 681 19 683 21
rect 718 20 720 22
rect 728 28 730 30
rect 752 35 754 37
rect 770 35 772 37
rect 793 27 795 29
rect 762 19 764 21
rect 781 19 783 21
rect 1 -40 3 -38
rect -10 -48 -8 -46
rect 11 -48 13 -46
rect 35 -55 37 -53
rect 45 -39 47 -37
rect 64 -39 66 -37
rect 53 -55 55 -53
rect 107 -40 109 -38
rect 76 -47 78 -45
rect 96 -48 98 -46
rect 117 -48 119 -46
rect 141 -55 143 -53
rect 151 -39 153 -37
rect 170 -39 172 -37
rect 159 -55 161 -53
rect 213 -40 215 -38
rect 182 -47 184 -45
rect 202 -48 204 -46
rect 223 -48 225 -46
rect 247 -55 249 -53
rect 257 -39 259 -37
rect 276 -39 278 -37
rect 265 -55 267 -53
rect 319 -40 321 -38
rect 288 -47 290 -45
rect 308 -48 310 -46
rect 329 -48 331 -46
rect 353 -55 355 -53
rect 363 -39 365 -37
rect 382 -39 384 -37
rect 371 -55 373 -53
rect 425 -40 427 -38
rect 394 -47 396 -45
rect 414 -48 416 -46
rect 435 -48 437 -46
rect 459 -55 461 -53
rect 469 -39 471 -37
rect 488 -39 490 -37
rect 477 -55 479 -53
rect 531 -40 533 -38
rect 500 -47 502 -45
rect 520 -48 522 -46
rect 541 -48 543 -46
rect 565 -55 567 -53
rect 575 -39 577 -37
rect 594 -39 596 -37
rect 583 -55 585 -53
rect 637 -40 639 -38
rect 606 -47 608 -45
rect 626 -48 628 -46
rect 647 -48 649 -46
rect 671 -55 673 -53
rect 681 -39 683 -37
rect 700 -39 702 -37
rect 689 -55 691 -53
rect 743 -40 745 -38
rect 712 -47 714 -45
rect 732 -48 734 -46
rect 753 -48 755 -46
rect 777 -55 779 -53
rect 787 -39 789 -37
rect 806 -39 808 -37
rect 795 -55 797 -53
rect 849 -40 851 -38
rect 818 -47 820 -45
rect 838 -48 840 -46
rect 859 -48 861 -46
rect 883 -55 885 -53
rect 893 -39 895 -37
rect 912 -39 914 -37
rect 901 -55 903 -53
rect 924 -47 926 -45
<< pdifct1 >>
rect 126 1138 128 1140
rect 153 1138 155 1140
rect 153 1131 155 1133
rect 186 1145 188 1147
rect 186 1138 188 1140
rect 274 1138 276 1140
rect 360 1146 362 1148
rect 310 1138 312 1140
rect 330 1138 332 1140
rect 330 1131 332 1133
rect 360 1139 362 1141
rect 341 1121 343 1123
rect 579 1139 581 1141
rect 650 1138 652 1140
rect 677 1146 679 1148
rect 677 1139 679 1141
rect 722 1145 724 1147
rect 722 1138 724 1140
rect 221 1109 223 1111
rect 118 1091 120 1093
rect 118 1084 120 1086
rect 146 1092 148 1094
rect 146 1085 148 1087
rect 261 1109 263 1111
rect 190 1093 192 1095
rect 190 1086 192 1088
rect 293 1091 295 1093
rect 585 1091 587 1093
rect 585 1084 587 1086
rect 603 1092 605 1094
rect 603 1085 605 1087
rect 695 1092 697 1094
rect 126 994 128 996
rect 218 994 220 996
rect 304 1000 306 1002
rect 304 993 306 995
rect 513 1002 515 1004
rect 513 995 515 997
rect 273 977 275 979
rect 598 1001 600 1003
rect 598 994 600 996
rect 659 1001 661 1003
rect 659 994 661 996
rect 675 1002 677 1004
rect 675 995 677 997
rect 722 1001 724 1003
rect 722 994 724 996
rect 85 955 87 957
rect 85 948 87 950
rect 118 947 120 949
rect 118 940 120 942
rect 146 948 148 950
rect 146 941 148 943
rect 212 948 214 950
rect 300 948 302 950
rect 300 941 302 943
rect 523 948 525 950
rect 581 948 583 950
rect 581 941 583 943
rect 636 948 638 950
rect 636 941 638 943
rect 656 948 658 950
rect 656 941 658 943
rect 695 948 697 950
rect 118 857 120 859
rect 118 850 120 852
rect 167 857 169 859
rect 167 850 169 852
rect 250 857 252 859
rect 250 850 252 852
rect 266 858 268 860
rect 266 851 268 853
rect 294 857 296 859
rect 294 850 296 852
rect 338 856 340 858
rect 338 849 340 851
rect 518 857 520 859
rect 518 850 520 852
rect 533 858 535 860
rect 533 851 535 853
rect 369 833 371 835
rect 591 857 593 859
rect 591 850 593 852
rect 609 857 611 859
rect 609 850 611 852
rect 695 856 697 858
rect 695 849 697 851
rect 664 833 666 835
rect 719 850 721 852
rect 719 843 721 845
rect 739 850 741 852
rect 739 843 741 845
rect 82 811 84 813
rect 82 804 84 806
rect 102 811 104 813
rect 102 804 104 806
rect 157 821 159 823
rect 126 805 128 807
rect 126 798 128 800
rect 212 804 214 806
rect 212 797 214 799
rect 230 804 232 806
rect 230 797 232 799
rect 452 821 454 823
rect 288 803 290 805
rect 288 796 290 798
rect 303 804 305 806
rect 303 797 305 799
rect 483 805 485 807
rect 483 798 485 800
rect 527 804 529 806
rect 527 797 529 799
rect 555 803 557 805
rect 555 796 557 798
rect 571 804 573 806
rect 571 797 573 799
rect 654 804 656 806
rect 654 797 656 799
rect 703 804 705 806
rect 703 797 705 799
rect 126 706 128 708
rect 165 713 167 715
rect 165 706 167 708
rect 185 713 187 715
rect 185 706 187 708
rect 240 713 242 715
rect 240 706 242 708
rect 298 706 300 708
rect 322 714 324 716
rect 322 707 324 709
rect 521 713 523 715
rect 521 706 523 708
rect 609 706 611 708
rect 675 713 677 715
rect 675 706 677 708
rect 703 714 705 716
rect 703 707 705 709
rect 736 706 738 708
rect 736 699 738 701
rect 99 660 101 662
rect 99 653 101 655
rect 146 659 148 661
rect 146 652 148 654
rect 162 660 164 662
rect 162 653 164 655
rect 223 660 225 662
rect 223 653 225 655
rect 548 677 550 679
rect 517 661 519 663
rect 517 654 519 656
rect 603 660 605 662
rect 695 660 697 662
rect 126 562 128 564
rect 218 569 220 571
rect 218 562 220 564
rect 236 570 238 572
rect 236 563 238 565
rect 528 563 530 565
rect 631 568 633 570
rect 631 561 633 563
rect 560 545 562 547
rect 675 569 677 571
rect 675 562 677 564
rect 703 570 705 572
rect 703 563 705 565
rect 600 545 602 547
rect 99 516 101 518
rect 99 509 101 511
rect 144 515 146 517
rect 144 508 146 510
rect 171 516 173 518
rect 242 515 244 517
rect 480 533 482 535
rect 461 515 463 517
rect 491 523 493 525
rect 491 516 493 518
rect 511 516 513 518
rect 461 508 463 510
rect 547 516 549 518
rect 635 516 637 518
rect 635 509 637 511
rect 668 523 670 525
rect 668 516 670 518
rect 695 516 697 518
rect 38 323 40 325
rect 38 316 40 318
rect 38 309 40 311
rect 107 316 109 318
rect 138 323 140 325
rect 138 316 140 318
rect 138 309 140 311
rect 238 323 240 325
rect 238 316 240 318
rect 238 309 240 311
rect 338 316 340 318
rect 338 309 340 311
rect 438 323 440 325
rect 438 316 440 318
rect 438 309 440 311
rect 538 323 540 325
rect 538 316 540 318
rect 538 309 540 311
rect 638 323 640 325
rect 638 316 640 318
rect 638 309 640 311
rect 738 323 740 325
rect 738 316 740 318
rect 738 309 740 311
rect 62 275 64 277
rect 62 268 64 270
rect 62 261 64 263
rect 162 275 164 277
rect 162 268 164 270
rect 162 261 164 263
rect 262 275 264 277
rect 262 268 264 270
rect 262 261 264 263
rect 362 275 364 277
rect 362 268 364 270
rect 362 261 364 263
rect 464 275 466 277
rect 464 268 466 270
rect 464 261 466 263
rect 564 275 566 277
rect 564 268 566 270
rect 564 261 566 263
rect 664 275 666 277
rect 664 268 666 270
rect 664 261 666 263
rect 764 275 766 277
rect 764 268 766 270
rect 764 261 766 263
rect 62 179 64 181
rect 62 172 64 174
rect 62 165 64 167
rect 162 179 164 181
rect 162 172 164 174
rect 162 165 164 167
rect 262 179 264 181
rect 262 172 264 174
rect 262 165 264 167
rect 362 179 364 181
rect 362 172 364 174
rect 362 165 364 167
rect 464 179 466 181
rect 464 172 466 174
rect 464 165 466 167
rect 564 179 566 181
rect 564 172 566 174
rect 564 165 566 167
rect 664 179 666 181
rect 664 172 666 174
rect 664 165 666 167
rect 764 179 766 181
rect 764 172 766 174
rect 764 165 766 167
rect 62 131 64 133
rect 62 124 64 126
rect 62 117 64 119
rect 162 131 164 133
rect 162 124 164 126
rect 162 117 164 119
rect 262 131 264 133
rect 262 124 264 126
rect 262 117 264 119
rect 362 131 364 133
rect 362 124 364 126
rect 362 117 364 119
rect 464 131 466 133
rect 464 124 466 126
rect 464 117 466 119
rect 564 131 566 133
rect 564 124 566 126
rect 564 117 566 119
rect 664 131 666 133
rect 664 124 666 126
rect 664 117 666 119
rect 764 131 766 133
rect 764 124 766 126
rect 764 117 766 119
rect 38 35 40 37
rect 38 28 40 30
rect 38 21 40 23
rect 107 28 109 30
rect 138 35 140 37
rect 138 28 140 30
rect 138 21 140 23
rect 238 35 240 37
rect 238 28 240 30
rect 238 21 240 23
rect 338 35 340 37
rect 338 28 340 30
rect 338 21 340 23
rect 438 35 440 37
rect 438 28 440 30
rect 438 21 440 23
rect 538 35 540 37
rect 538 28 540 30
rect 538 21 540 23
rect 638 35 640 37
rect 638 28 640 30
rect 638 21 640 23
rect 738 35 740 37
rect 738 28 740 30
rect 738 21 740 23
rect 21 -41 23 -39
rect 21 -48 23 -46
rect 21 -55 23 -53
rect 127 -41 129 -39
rect 127 -48 129 -46
rect 127 -55 129 -53
rect 233 -41 235 -39
rect 233 -48 235 -46
rect 233 -55 235 -53
rect 339 -41 341 -39
rect 339 -48 341 -46
rect 339 -55 341 -53
rect 445 -41 447 -39
rect 445 -48 447 -46
rect 445 -55 447 -53
rect 551 -41 553 -39
rect 551 -48 553 -46
rect 551 -55 553 -53
rect 657 -41 659 -39
rect 657 -48 659 -46
rect 657 -55 659 -53
rect 763 -41 765 -39
rect 763 -48 765 -46
rect 763 -55 765 -53
rect 869 -41 871 -39
rect 869 -48 871 -46
rect 869 -55 871 -53
<< alu0 >>
rect 94 1174 100 1180
rect 94 1172 96 1174
rect 98 1172 100 1174
rect 94 1171 100 1172
rect 107 1171 111 1173
rect 107 1169 108 1171
rect 110 1169 111 1171
rect 81 1166 85 1168
rect 81 1164 82 1166
rect 84 1164 85 1166
rect 81 1158 85 1164
rect 107 1166 111 1169
rect 107 1162 131 1166
rect 81 1154 92 1158
rect 88 1148 92 1154
rect 127 1158 131 1162
rect 107 1157 123 1158
rect 107 1155 119 1157
rect 121 1155 123 1157
rect 107 1154 123 1155
rect 127 1156 132 1158
rect 127 1154 129 1156
rect 131 1154 132 1156
rect 107 1148 111 1154
rect 127 1152 132 1154
rect 127 1150 131 1152
rect 88 1147 111 1148
rect 88 1145 90 1147
rect 92 1145 111 1147
rect 88 1144 111 1145
rect 99 1133 103 1135
rect 99 1131 100 1133
rect 102 1131 103 1133
rect 99 1126 103 1131
rect 107 1133 111 1144
rect 115 1147 131 1150
rect 115 1145 116 1147
rect 118 1146 131 1147
rect 118 1145 119 1146
rect 115 1140 119 1145
rect 115 1138 116 1140
rect 118 1138 119 1140
rect 115 1136 119 1138
rect 171 1171 175 1180
rect 171 1169 172 1171
rect 174 1169 175 1171
rect 171 1167 175 1169
rect 242 1174 248 1180
rect 200 1173 220 1174
rect 200 1171 216 1173
rect 218 1171 220 1173
rect 242 1172 244 1174
rect 246 1172 248 1174
rect 242 1171 248 1172
rect 255 1171 259 1173
rect 200 1170 220 1171
rect 188 1167 189 1169
rect 200 1166 204 1170
rect 255 1169 256 1171
rect 258 1169 259 1171
rect 192 1162 204 1166
rect 192 1157 196 1162
rect 192 1155 193 1157
rect 195 1155 196 1157
rect 192 1143 196 1155
rect 229 1166 233 1168
rect 229 1164 230 1166
rect 232 1164 233 1166
rect 229 1158 233 1164
rect 255 1166 259 1169
rect 255 1162 279 1166
rect 229 1154 240 1158
rect 192 1140 209 1143
rect 192 1139 206 1140
rect 205 1138 206 1139
rect 208 1138 209 1140
rect 194 1135 200 1136
rect 107 1132 140 1133
rect 107 1130 136 1132
rect 138 1130 140 1132
rect 171 1133 175 1135
rect 171 1131 172 1133
rect 174 1131 175 1133
rect 107 1129 140 1130
rect 99 1124 100 1126
rect 102 1124 103 1126
rect 171 1126 175 1131
rect 171 1124 172 1126
rect 174 1124 175 1126
rect 194 1133 196 1135
rect 198 1133 200 1135
rect 194 1124 200 1133
rect 205 1133 209 1138
rect 236 1148 240 1154
rect 275 1158 279 1162
rect 255 1157 271 1158
rect 255 1155 267 1157
rect 269 1155 271 1157
rect 255 1154 271 1155
rect 275 1156 280 1158
rect 275 1154 277 1156
rect 279 1154 280 1156
rect 255 1148 259 1154
rect 275 1152 280 1154
rect 275 1150 279 1152
rect 236 1147 259 1148
rect 236 1145 238 1147
rect 240 1145 259 1147
rect 236 1144 259 1145
rect 205 1131 206 1133
rect 208 1131 209 1133
rect 205 1129 209 1131
rect 214 1133 220 1134
rect 214 1131 216 1133
rect 218 1131 220 1133
rect 214 1124 220 1131
rect 247 1133 251 1135
rect 247 1131 248 1133
rect 250 1131 251 1133
rect 247 1126 251 1131
rect 255 1133 259 1144
rect 263 1147 279 1150
rect 263 1145 264 1147
rect 266 1146 279 1147
rect 266 1145 267 1146
rect 263 1140 267 1145
rect 263 1138 264 1140
rect 266 1138 267 1140
rect 263 1136 267 1138
rect 325 1150 330 1151
rect 325 1148 327 1150
rect 329 1148 330 1150
rect 373 1169 377 1180
rect 566 1173 572 1180
rect 566 1171 568 1173
rect 570 1171 572 1173
rect 566 1170 572 1171
rect 589 1170 593 1180
rect 618 1174 624 1180
rect 618 1172 620 1174
rect 622 1172 624 1174
rect 618 1171 624 1172
rect 631 1171 635 1173
rect 325 1147 330 1148
rect 309 1133 313 1137
rect 255 1132 288 1133
rect 255 1130 284 1132
rect 286 1130 288 1132
rect 255 1129 288 1130
rect 299 1130 303 1132
rect 247 1124 248 1126
rect 250 1124 251 1126
rect 299 1128 300 1130
rect 302 1128 303 1130
rect 309 1131 310 1133
rect 312 1131 313 1133
rect 309 1129 313 1131
rect 319 1130 323 1132
rect 299 1124 303 1128
rect 319 1128 320 1130
rect 322 1128 323 1130
rect 362 1162 363 1168
rect 373 1167 374 1169
rect 376 1167 377 1169
rect 589 1168 590 1170
rect 592 1168 593 1170
rect 631 1169 632 1171
rect 634 1169 635 1171
rect 373 1165 377 1167
rect 589 1166 593 1168
rect 605 1166 609 1168
rect 605 1164 606 1166
rect 608 1164 609 1166
rect 362 1143 363 1150
rect 588 1150 590 1157
rect 605 1158 609 1164
rect 631 1166 635 1169
rect 631 1162 655 1166
rect 605 1154 616 1158
rect 587 1142 593 1143
rect 587 1140 589 1142
rect 591 1140 593 1142
rect 587 1135 593 1140
rect 567 1134 573 1135
rect 369 1133 375 1134
rect 369 1131 371 1133
rect 373 1131 375 1133
rect 319 1124 323 1128
rect 369 1124 375 1131
rect 567 1132 569 1134
rect 571 1132 573 1134
rect 567 1127 573 1132
rect 567 1125 569 1127
rect 571 1125 573 1127
rect 567 1124 573 1125
rect 587 1133 589 1135
rect 591 1133 593 1135
rect 587 1124 593 1133
rect 612 1148 616 1154
rect 651 1158 655 1162
rect 631 1157 647 1158
rect 631 1155 643 1157
rect 645 1155 647 1157
rect 631 1154 647 1155
rect 651 1156 656 1158
rect 651 1154 653 1156
rect 655 1154 656 1156
rect 631 1148 635 1154
rect 651 1152 656 1154
rect 651 1150 655 1152
rect 612 1147 635 1148
rect 612 1145 614 1147
rect 616 1145 635 1147
rect 612 1144 635 1145
rect 623 1133 627 1135
rect 623 1131 624 1133
rect 626 1131 627 1133
rect 623 1126 627 1131
rect 631 1133 635 1144
rect 639 1147 655 1150
rect 639 1145 640 1147
rect 642 1146 655 1147
rect 642 1145 643 1146
rect 639 1140 643 1145
rect 639 1138 640 1140
rect 642 1138 643 1140
rect 639 1136 643 1138
rect 690 1169 694 1180
rect 715 1178 717 1180
rect 719 1178 721 1180
rect 679 1162 680 1168
rect 690 1167 691 1169
rect 693 1167 694 1169
rect 690 1165 694 1167
rect 715 1173 721 1178
rect 735 1178 737 1180
rect 739 1178 741 1180
rect 735 1177 741 1178
rect 715 1171 717 1173
rect 719 1171 721 1173
rect 715 1170 721 1171
rect 679 1143 680 1150
rect 686 1133 692 1134
rect 631 1132 664 1133
rect 631 1130 660 1132
rect 662 1130 664 1132
rect 631 1129 664 1130
rect 686 1131 688 1133
rect 690 1131 692 1133
rect 623 1124 624 1126
rect 626 1124 627 1126
rect 686 1124 692 1131
rect 703 1133 709 1134
rect 703 1131 705 1133
rect 707 1131 709 1133
rect 703 1126 709 1131
rect 703 1124 705 1126
rect 707 1124 709 1126
rect 737 1133 743 1134
rect 737 1131 739 1133
rect 741 1131 743 1133
rect 737 1126 743 1131
rect 737 1124 739 1126
rect 741 1124 743 1126
rect 80 1106 82 1108
rect 84 1106 86 1108
rect 80 1101 86 1106
rect 100 1106 102 1108
rect 104 1106 106 1108
rect 80 1099 82 1101
rect 84 1099 86 1101
rect 80 1098 86 1099
rect 91 1101 95 1103
rect 91 1099 92 1101
rect 94 1099 95 1101
rect 91 1095 95 1099
rect 100 1101 106 1106
rect 100 1099 102 1101
rect 104 1099 106 1101
rect 100 1098 106 1099
rect 127 1101 133 1108
rect 127 1099 129 1101
rect 131 1099 133 1101
rect 127 1098 133 1099
rect 154 1099 160 1108
rect 154 1097 156 1099
rect 158 1097 160 1099
rect 154 1096 160 1097
rect 165 1101 169 1103
rect 165 1099 166 1101
rect 168 1099 169 1101
rect 92 1094 95 1095
rect 94 1092 95 1094
rect 92 1090 95 1092
rect 165 1094 169 1099
rect 174 1101 180 1108
rect 174 1099 176 1101
rect 178 1099 180 1101
rect 174 1098 180 1099
rect 198 1100 204 1108
rect 198 1098 200 1100
rect 202 1098 204 1100
rect 198 1097 204 1098
rect 209 1100 236 1102
rect 209 1098 210 1100
rect 212 1099 236 1100
rect 212 1098 232 1099
rect 165 1093 166 1094
rect 103 1077 104 1081
rect 120 1082 121 1089
rect 152 1092 166 1093
rect 168 1092 169 1094
rect 152 1089 169 1092
rect 103 1061 107 1063
rect 103 1059 104 1061
rect 106 1059 107 1061
rect 103 1054 107 1059
rect 120 1064 121 1070
rect 131 1065 135 1067
rect 131 1063 132 1065
rect 134 1063 135 1065
rect 103 1052 104 1054
rect 106 1052 107 1054
rect 131 1052 135 1063
rect 152 1077 156 1089
rect 209 1093 213 1098
rect 230 1097 232 1098
rect 234 1097 236 1099
rect 204 1091 210 1093
rect 212 1091 213 1093
rect 152 1075 153 1077
rect 155 1075 156 1077
rect 152 1070 156 1075
rect 152 1066 164 1070
rect 148 1063 149 1065
rect 160 1062 164 1066
rect 192 1084 193 1090
rect 204 1089 213 1091
rect 204 1086 208 1089
rect 230 1092 236 1097
rect 230 1090 232 1092
rect 234 1090 236 1092
rect 230 1089 236 1090
rect 196 1082 208 1086
rect 196 1077 200 1082
rect 215 1081 221 1082
rect 196 1075 197 1077
rect 199 1075 200 1077
rect 196 1069 200 1075
rect 160 1061 180 1062
rect 160 1059 176 1061
rect 178 1059 180 1061
rect 160 1058 180 1059
rect 192 1063 193 1069
rect 196 1065 205 1069
rect 260 1074 261 1080
rect 201 1061 205 1065
rect 322 1099 328 1108
rect 322 1097 324 1099
rect 326 1097 328 1099
rect 572 1101 578 1108
rect 572 1099 574 1101
rect 576 1099 578 1101
rect 572 1098 578 1099
rect 611 1099 617 1108
rect 322 1092 328 1097
rect 611 1097 613 1099
rect 615 1097 617 1099
rect 611 1096 617 1097
rect 622 1101 626 1103
rect 622 1099 623 1101
rect 625 1099 626 1101
rect 322 1090 324 1092
rect 326 1090 328 1092
rect 322 1089 328 1090
rect 584 1082 585 1089
rect 201 1060 231 1061
rect 201 1058 227 1060
rect 229 1058 231 1060
rect 201 1057 231 1058
rect 257 1060 261 1062
rect 257 1058 258 1060
rect 260 1058 261 1060
rect 257 1052 261 1058
rect 299 1060 303 1062
rect 299 1058 300 1060
rect 302 1058 303 1060
rect 299 1052 303 1058
rect 570 1065 574 1067
rect 570 1063 571 1065
rect 573 1063 574 1065
rect 584 1064 585 1070
rect 570 1052 574 1063
rect 622 1094 626 1099
rect 631 1101 637 1108
rect 631 1099 633 1101
rect 635 1099 637 1101
rect 631 1098 637 1099
rect 649 1106 651 1108
rect 653 1106 655 1108
rect 649 1101 655 1106
rect 669 1106 671 1108
rect 673 1106 675 1108
rect 649 1099 651 1101
rect 653 1099 655 1101
rect 649 1098 655 1099
rect 660 1101 664 1103
rect 660 1099 661 1101
rect 663 1099 664 1101
rect 660 1095 664 1099
rect 669 1101 675 1106
rect 720 1106 721 1108
rect 723 1106 724 1108
rect 669 1099 671 1101
rect 673 1099 675 1101
rect 683 1102 716 1103
rect 683 1100 685 1102
rect 687 1100 716 1102
rect 683 1099 716 1100
rect 669 1098 675 1099
rect 622 1093 623 1094
rect 609 1092 623 1093
rect 625 1092 626 1094
rect 609 1089 626 1092
rect 609 1077 613 1089
rect 660 1094 663 1095
rect 660 1092 661 1094
rect 660 1090 663 1092
rect 609 1075 610 1077
rect 612 1075 613 1077
rect 609 1070 613 1075
rect 609 1066 621 1070
rect 605 1063 606 1065
rect 617 1062 621 1066
rect 651 1077 652 1081
rect 617 1061 637 1062
rect 617 1059 633 1061
rect 635 1059 637 1061
rect 617 1058 637 1059
rect 648 1061 652 1063
rect 648 1059 649 1061
rect 651 1059 652 1061
rect 648 1054 652 1059
rect 704 1094 708 1096
rect 704 1092 705 1094
rect 707 1092 708 1094
rect 704 1087 708 1092
rect 704 1086 705 1087
rect 692 1085 705 1086
rect 707 1085 708 1087
rect 692 1082 708 1085
rect 712 1088 716 1099
rect 720 1101 724 1106
rect 720 1099 721 1101
rect 723 1099 724 1101
rect 720 1097 724 1099
rect 712 1087 735 1088
rect 712 1085 731 1087
rect 733 1085 735 1087
rect 712 1084 735 1085
rect 692 1080 696 1082
rect 691 1078 696 1080
rect 712 1078 716 1084
rect 691 1076 692 1078
rect 694 1076 696 1078
rect 691 1074 696 1076
rect 700 1077 716 1078
rect 700 1075 702 1077
rect 704 1075 716 1077
rect 700 1074 716 1075
rect 692 1070 696 1074
rect 731 1078 735 1084
rect 731 1074 742 1078
rect 692 1066 716 1070
rect 712 1063 716 1066
rect 738 1068 742 1074
rect 738 1066 739 1068
rect 741 1066 742 1068
rect 738 1064 742 1066
rect 712 1061 713 1063
rect 715 1061 716 1063
rect 712 1059 716 1061
rect 723 1060 729 1061
rect 723 1058 725 1060
rect 727 1058 729 1060
rect 648 1052 649 1054
rect 651 1052 652 1054
rect 723 1052 729 1058
rect 94 1030 100 1036
rect 171 1034 172 1036
rect 174 1034 175 1036
rect 94 1028 96 1030
rect 98 1028 100 1030
rect 94 1027 100 1028
rect 107 1027 111 1029
rect 107 1025 108 1027
rect 110 1025 111 1027
rect 81 1022 85 1024
rect 81 1020 82 1022
rect 84 1020 85 1022
rect 81 1014 85 1020
rect 107 1022 111 1025
rect 107 1018 131 1022
rect 81 1010 92 1014
rect 88 1004 92 1010
rect 127 1014 131 1018
rect 107 1013 123 1014
rect 107 1011 119 1013
rect 121 1011 123 1013
rect 107 1010 123 1011
rect 127 1012 132 1014
rect 127 1010 129 1012
rect 131 1010 132 1012
rect 107 1004 111 1010
rect 127 1008 132 1010
rect 127 1006 131 1008
rect 88 1003 111 1004
rect 88 1001 90 1003
rect 92 1001 111 1003
rect 88 1000 111 1001
rect 99 989 103 991
rect 99 987 100 989
rect 102 987 103 989
rect 99 982 103 987
rect 107 989 111 1000
rect 115 1003 131 1006
rect 115 1001 116 1003
rect 118 1002 131 1003
rect 118 1001 119 1002
rect 115 996 119 1001
rect 115 994 116 996
rect 118 994 119 996
rect 115 992 119 994
rect 171 1029 175 1034
rect 171 1027 172 1029
rect 174 1027 175 1029
rect 171 1025 175 1027
rect 265 1030 295 1031
rect 265 1028 267 1030
rect 269 1028 295 1030
rect 265 1027 295 1028
rect 171 1007 172 1011
rect 291 1023 295 1027
rect 291 1019 300 1023
rect 303 1019 304 1025
rect 296 1013 300 1019
rect 296 1011 297 1013
rect 299 1011 300 1013
rect 275 1006 281 1007
rect 296 1006 300 1011
rect 288 1002 300 1006
rect 160 996 163 998
rect 162 994 163 996
rect 260 998 266 999
rect 260 996 262 998
rect 264 996 266 998
rect 160 993 163 994
rect 148 989 154 990
rect 107 988 140 989
rect 107 986 136 988
rect 138 986 140 988
rect 107 985 140 986
rect 148 987 150 989
rect 152 987 154 989
rect 99 980 100 982
rect 102 980 103 982
rect 148 982 154 987
rect 159 989 163 993
rect 159 987 160 989
rect 162 987 163 989
rect 159 985 163 987
rect 168 989 174 990
rect 168 987 170 989
rect 172 987 174 989
rect 148 980 150 982
rect 152 980 154 982
rect 168 982 174 987
rect 168 980 170 982
rect 172 980 174 982
rect 192 989 198 990
rect 192 987 194 989
rect 196 987 198 989
rect 192 982 198 987
rect 217 989 221 994
rect 260 991 266 996
rect 288 999 292 1002
rect 283 997 292 999
rect 303 998 304 1004
rect 283 995 284 997
rect 286 995 292 997
rect 217 987 218 989
rect 220 987 221 989
rect 217 985 221 987
rect 240 989 246 990
rect 240 987 242 989
rect 244 987 246 989
rect 192 980 194 982
rect 196 980 198 982
rect 240 982 246 987
rect 260 989 262 991
rect 264 990 266 991
rect 283 990 287 995
rect 526 1025 530 1036
rect 591 1034 593 1036
rect 595 1034 597 1036
rect 515 1018 516 1024
rect 526 1023 527 1025
rect 529 1023 530 1025
rect 526 1021 530 1023
rect 591 1029 597 1034
rect 611 1034 613 1036
rect 615 1034 617 1036
rect 611 1033 617 1034
rect 591 1027 593 1029
rect 595 1027 597 1029
rect 591 1026 597 1027
rect 627 1029 647 1030
rect 627 1027 629 1029
rect 631 1027 647 1029
rect 627 1026 647 1027
rect 515 999 516 1006
rect 643 1022 647 1026
rect 658 1023 659 1025
rect 643 1018 655 1022
rect 651 1013 655 1018
rect 651 1011 652 1013
rect 654 1011 655 1013
rect 264 989 284 990
rect 260 988 284 989
rect 286 988 287 990
rect 260 986 287 988
rect 292 990 298 991
rect 292 988 294 990
rect 296 988 298 990
rect 240 980 242 982
rect 244 980 246 982
rect 292 980 298 988
rect 651 999 655 1011
rect 638 996 655 999
rect 638 994 639 996
rect 641 995 655 996
rect 688 1025 692 1036
rect 715 1034 717 1036
rect 719 1034 721 1036
rect 677 1018 678 1024
rect 688 1023 689 1025
rect 691 1023 692 1025
rect 688 1021 692 1023
rect 715 1029 721 1034
rect 735 1034 737 1036
rect 739 1034 741 1036
rect 735 1033 741 1034
rect 715 1027 717 1029
rect 719 1027 721 1029
rect 715 1026 721 1027
rect 677 999 678 1006
rect 641 994 642 995
rect 522 989 528 990
rect 522 987 524 989
rect 526 987 528 989
rect 522 980 528 987
rect 579 989 585 990
rect 579 987 581 989
rect 583 987 585 989
rect 579 982 585 987
rect 579 980 581 982
rect 583 980 585 982
rect 613 989 619 990
rect 613 987 615 989
rect 617 987 619 989
rect 613 982 619 987
rect 613 980 615 982
rect 617 980 619 982
rect 627 989 633 990
rect 627 987 629 989
rect 631 987 633 989
rect 627 980 633 987
rect 638 989 642 994
rect 638 987 639 989
rect 641 987 642 989
rect 638 985 642 987
rect 647 991 653 992
rect 647 989 649 991
rect 651 989 653 991
rect 647 980 653 989
rect 684 989 690 990
rect 684 987 686 989
rect 688 987 690 989
rect 684 980 690 987
rect 703 989 709 990
rect 703 987 705 989
rect 707 987 709 989
rect 703 982 709 987
rect 703 980 705 982
rect 707 980 709 982
rect 737 989 743 990
rect 737 987 739 989
rect 741 987 743 989
rect 737 982 743 987
rect 737 980 739 982
rect 741 980 743 982
rect 103 962 104 964
rect 106 962 107 964
rect 103 957 107 962
rect 103 955 104 957
rect 106 955 107 957
rect 103 953 107 955
rect 127 957 133 964
rect 127 955 129 957
rect 131 955 133 957
rect 127 954 133 955
rect 154 955 160 964
rect 154 953 156 955
rect 158 953 160 955
rect 154 952 160 953
rect 165 957 169 959
rect 165 955 166 957
rect 168 955 169 957
rect 165 950 169 955
rect 174 957 180 964
rect 237 962 238 964
rect 240 962 241 964
rect 174 955 176 957
rect 178 955 180 957
rect 200 958 233 959
rect 200 956 202 958
rect 204 956 233 958
rect 200 955 233 956
rect 174 954 180 955
rect 165 949 166 950
rect 120 938 121 945
rect 152 948 166 949
rect 168 948 169 950
rect 152 945 169 948
rect 103 919 107 921
rect 103 917 104 919
rect 106 917 107 919
rect 103 908 107 917
rect 120 920 121 926
rect 131 921 135 923
rect 131 919 132 921
rect 134 919 135 921
rect 131 908 135 919
rect 152 933 156 945
rect 221 950 225 952
rect 221 948 222 950
rect 224 948 225 950
rect 221 943 225 948
rect 221 942 222 943
rect 209 941 222 942
rect 224 941 225 943
rect 209 938 225 941
rect 229 944 233 955
rect 237 957 241 962
rect 237 955 238 957
rect 240 955 241 957
rect 237 953 241 955
rect 268 957 274 964
rect 268 955 270 957
rect 272 955 274 957
rect 268 954 274 955
rect 279 957 283 959
rect 279 955 280 957
rect 282 955 283 957
rect 229 943 252 944
rect 229 941 248 943
rect 250 941 252 943
rect 229 940 252 941
rect 209 936 213 938
rect 152 931 153 933
rect 155 931 156 933
rect 152 926 156 931
rect 152 922 164 926
rect 148 919 149 921
rect 160 918 164 922
rect 160 917 180 918
rect 160 915 176 917
rect 178 915 180 917
rect 160 914 180 915
rect 208 934 213 936
rect 229 934 233 940
rect 208 932 209 934
rect 211 932 213 934
rect 208 930 213 932
rect 217 933 233 934
rect 217 931 219 933
rect 221 931 233 933
rect 217 930 233 931
rect 209 926 213 930
rect 248 934 252 940
rect 279 950 283 955
rect 288 955 294 964
rect 548 962 549 964
rect 551 962 552 964
rect 511 958 544 959
rect 511 956 513 958
rect 515 956 544 958
rect 511 955 544 956
rect 288 953 290 955
rect 292 953 294 955
rect 288 952 294 953
rect 279 948 280 950
rect 282 949 283 950
rect 282 948 296 949
rect 279 945 296 948
rect 248 930 259 934
rect 209 922 233 926
rect 229 919 233 922
rect 255 924 259 930
rect 255 922 256 924
rect 258 922 259 924
rect 255 920 259 922
rect 292 933 296 945
rect 292 931 293 933
rect 295 931 296 933
rect 292 926 296 931
rect 284 922 296 926
rect 229 917 230 919
rect 232 917 233 919
rect 284 918 288 922
rect 299 919 300 921
rect 268 917 288 918
rect 229 915 233 917
rect 240 916 246 917
rect 240 914 242 916
rect 244 914 246 916
rect 268 915 270 917
rect 272 915 288 917
rect 268 914 288 915
rect 240 908 246 914
rect 532 950 536 952
rect 532 948 533 950
rect 535 948 536 950
rect 532 943 536 948
rect 532 942 533 943
rect 520 941 533 942
rect 535 941 536 943
rect 520 938 536 941
rect 540 944 544 955
rect 548 957 552 962
rect 548 955 549 957
rect 551 955 552 957
rect 548 953 552 955
rect 540 943 563 944
rect 540 941 559 943
rect 561 941 563 943
rect 540 940 563 941
rect 520 936 524 938
rect 519 934 524 936
rect 540 934 544 940
rect 519 932 520 934
rect 522 932 524 934
rect 519 930 524 932
rect 528 933 544 934
rect 528 931 530 933
rect 532 931 544 933
rect 528 930 544 931
rect 520 926 524 930
rect 559 934 563 940
rect 589 955 595 964
rect 589 953 591 955
rect 593 953 595 955
rect 589 952 595 953
rect 600 957 604 959
rect 600 955 601 957
rect 603 955 604 957
rect 600 950 604 955
rect 609 957 615 964
rect 609 955 611 957
rect 613 955 615 957
rect 609 954 615 955
rect 625 955 629 964
rect 625 953 626 955
rect 628 953 629 955
rect 625 951 629 953
rect 644 955 650 964
rect 644 953 646 955
rect 648 953 650 955
rect 600 949 601 950
rect 587 948 601 949
rect 603 948 604 950
rect 587 945 604 948
rect 559 930 570 934
rect 520 922 544 926
rect 540 919 544 922
rect 566 924 570 930
rect 566 922 567 924
rect 569 922 570 924
rect 566 920 570 922
rect 540 917 541 919
rect 543 917 544 919
rect 587 933 591 945
rect 644 948 650 953
rect 665 955 669 964
rect 720 962 721 964
rect 723 962 724 964
rect 683 958 716 959
rect 683 956 685 958
rect 687 956 716 958
rect 683 955 716 956
rect 665 953 666 955
rect 668 953 669 955
rect 644 946 646 948
rect 648 946 650 948
rect 644 945 650 946
rect 665 948 669 953
rect 665 946 666 948
rect 668 946 669 948
rect 665 944 669 946
rect 704 950 708 952
rect 704 948 705 950
rect 707 948 708 950
rect 587 931 588 933
rect 590 931 591 933
rect 587 926 591 931
rect 587 922 599 926
rect 583 919 584 921
rect 540 915 544 917
rect 551 916 557 917
rect 551 914 553 916
rect 555 914 557 916
rect 551 908 557 914
rect 595 918 599 922
rect 623 924 649 925
rect 623 922 625 924
rect 627 923 649 924
rect 627 922 646 923
rect 623 921 646 922
rect 648 921 649 923
rect 595 917 615 918
rect 644 917 649 921
rect 704 943 708 948
rect 704 942 705 943
rect 692 941 705 942
rect 707 941 708 943
rect 692 938 708 941
rect 712 944 716 955
rect 720 957 724 962
rect 720 955 721 957
rect 723 955 724 957
rect 720 953 724 955
rect 712 943 735 944
rect 712 941 731 943
rect 733 941 735 943
rect 712 940 735 941
rect 692 936 696 938
rect 691 934 696 936
rect 712 934 716 940
rect 691 932 692 934
rect 694 932 696 934
rect 691 930 696 932
rect 700 933 716 934
rect 700 931 702 933
rect 704 931 716 933
rect 700 930 716 931
rect 692 926 696 930
rect 731 934 735 940
rect 731 930 742 934
rect 692 922 716 926
rect 712 919 716 922
rect 738 924 742 930
rect 738 922 739 924
rect 741 922 742 924
rect 738 920 742 922
rect 595 915 611 917
rect 613 915 615 917
rect 595 914 615 915
rect 635 915 639 917
rect 635 913 636 915
rect 638 913 639 915
rect 644 916 670 917
rect 644 914 646 916
rect 648 914 666 916
rect 668 914 670 916
rect 712 917 713 919
rect 715 917 716 919
rect 712 915 716 917
rect 723 916 729 917
rect 723 914 725 916
rect 727 914 729 916
rect 644 913 670 914
rect 635 908 639 913
rect 723 908 729 914
rect 82 891 86 892
rect 82 889 83 891
rect 85 889 86 891
rect 82 887 86 889
rect 81 854 87 855
rect 81 852 83 854
rect 85 852 87 854
rect 81 847 87 852
rect 81 845 83 847
rect 85 845 87 847
rect 81 836 87 845
rect 92 854 105 855
rect 92 852 94 854
rect 92 850 96 852
rect 132 885 152 886
rect 132 883 148 885
rect 150 883 152 885
rect 132 882 152 883
rect 120 879 121 881
rect 132 878 136 882
rect 181 885 201 886
rect 181 883 197 885
rect 199 883 201 885
rect 181 882 201 883
rect 218 885 238 886
rect 218 883 220 885
rect 222 883 238 885
rect 218 882 238 883
rect 124 874 136 878
rect 124 869 128 874
rect 124 867 125 869
rect 127 867 128 869
rect 124 855 128 867
rect 124 852 141 855
rect 124 851 138 852
rect 92 847 98 850
rect 92 845 94 847
rect 96 845 98 847
rect 137 850 138 851
rect 140 850 141 852
rect 92 844 98 845
rect 103 845 109 846
rect 103 843 105 845
rect 107 843 109 845
rect 126 847 132 848
rect 126 845 128 847
rect 130 845 132 847
rect 103 836 109 843
rect 126 836 132 845
rect 137 845 141 850
rect 169 879 170 881
rect 181 878 185 882
rect 173 874 185 878
rect 173 869 177 874
rect 173 867 174 869
rect 176 867 177 869
rect 173 855 177 867
rect 234 878 238 882
rect 249 879 250 881
rect 234 874 246 878
rect 242 869 246 874
rect 242 867 243 869
rect 245 867 246 869
rect 173 852 190 855
rect 173 851 187 852
rect 186 850 187 851
rect 189 850 190 852
rect 175 847 181 848
rect 137 843 138 845
rect 140 843 141 845
rect 137 841 141 843
rect 146 845 152 846
rect 146 843 148 845
rect 150 843 152 845
rect 146 836 152 843
rect 175 845 177 847
rect 179 845 181 847
rect 175 836 181 845
rect 186 845 190 850
rect 242 855 246 867
rect 229 852 246 855
rect 229 850 230 852
rect 232 851 246 852
rect 232 850 233 851
rect 186 843 187 845
rect 189 843 190 845
rect 186 841 190 843
rect 195 845 201 846
rect 195 843 197 845
rect 199 843 201 845
rect 195 836 201 843
rect 218 845 224 846
rect 218 843 220 845
rect 222 843 224 845
rect 218 836 224 843
rect 229 845 233 850
rect 279 881 283 892
rect 268 874 269 880
rect 279 879 280 881
rect 282 879 283 881
rect 279 877 283 879
rect 308 885 328 886
rect 308 883 324 885
rect 326 883 328 885
rect 308 882 328 883
rect 268 855 269 862
rect 296 879 297 881
rect 308 878 312 882
rect 349 886 379 887
rect 349 884 375 886
rect 377 884 379 886
rect 349 883 379 884
rect 486 885 506 886
rect 486 883 488 885
rect 490 883 506 885
rect 300 874 312 878
rect 300 869 304 874
rect 300 867 301 869
rect 303 867 304 869
rect 300 855 304 867
rect 300 852 317 855
rect 300 851 314 852
rect 313 850 314 851
rect 316 850 317 852
rect 229 843 230 845
rect 232 843 233 845
rect 229 841 233 843
rect 238 847 244 848
rect 238 845 240 847
rect 242 845 244 847
rect 302 847 308 848
rect 238 836 244 845
rect 275 845 281 846
rect 275 843 277 845
rect 279 843 281 845
rect 275 836 281 843
rect 302 845 304 847
rect 306 845 308 847
rect 302 836 308 845
rect 313 845 317 850
rect 340 875 341 881
rect 349 879 353 883
rect 486 882 506 883
rect 344 875 353 879
rect 344 869 348 875
rect 344 867 345 869
rect 347 867 348 869
rect 344 862 348 867
rect 502 878 506 882
rect 517 879 518 881
rect 502 874 514 878
rect 510 869 514 874
rect 510 867 511 869
rect 513 867 514 869
rect 363 862 369 863
rect 340 854 341 860
rect 344 858 356 862
rect 352 855 356 858
rect 352 853 361 855
rect 352 851 358 853
rect 360 851 361 853
rect 313 843 314 845
rect 316 843 317 845
rect 313 841 317 843
rect 322 845 328 846
rect 322 843 324 845
rect 326 843 328 845
rect 322 836 328 843
rect 346 846 352 847
rect 346 844 348 846
rect 350 844 352 846
rect 346 836 352 844
rect 357 846 361 851
rect 378 854 384 855
rect 378 852 380 854
rect 382 852 384 854
rect 378 847 384 852
rect 510 855 514 867
rect 497 852 514 855
rect 497 850 498 852
rect 500 851 514 852
rect 500 850 501 851
rect 378 846 380 847
rect 357 844 358 846
rect 360 845 380 846
rect 382 845 384 847
rect 360 844 384 845
rect 357 842 384 844
rect 486 845 492 846
rect 486 843 488 845
rect 490 843 492 845
rect 486 836 492 843
rect 497 845 501 850
rect 546 881 550 892
rect 709 891 711 892
rect 713 891 715 892
rect 709 890 715 891
rect 559 885 579 886
rect 559 883 561 885
rect 563 883 579 885
rect 559 882 579 883
rect 535 874 536 880
rect 546 879 547 881
rect 549 879 550 881
rect 546 877 550 879
rect 575 878 579 882
rect 590 879 591 881
rect 575 874 587 878
rect 583 869 587 874
rect 583 867 584 869
rect 586 867 587 869
rect 535 855 536 862
rect 583 855 587 867
rect 570 852 587 855
rect 570 850 571 852
rect 573 851 587 852
rect 573 850 574 851
rect 497 843 498 845
rect 500 843 501 845
rect 497 841 501 843
rect 506 847 512 848
rect 506 845 508 847
rect 510 845 512 847
rect 506 836 512 845
rect 542 845 548 846
rect 542 843 544 845
rect 546 843 548 845
rect 542 836 548 843
rect 559 845 565 846
rect 559 843 561 845
rect 563 843 565 845
rect 559 836 565 843
rect 570 845 574 850
rect 656 886 686 887
rect 623 885 643 886
rect 623 883 639 885
rect 641 883 643 885
rect 656 884 658 886
rect 660 884 686 886
rect 656 883 686 884
rect 623 882 643 883
rect 611 879 612 881
rect 623 878 627 882
rect 682 879 686 883
rect 615 874 627 878
rect 615 869 619 874
rect 615 867 616 869
rect 618 867 619 869
rect 615 855 619 867
rect 682 875 691 879
rect 694 875 695 881
rect 687 869 691 875
rect 687 867 688 869
rect 690 867 691 869
rect 666 862 672 863
rect 687 862 691 867
rect 679 858 691 862
rect 615 852 632 855
rect 615 851 629 852
rect 628 850 629 851
rect 631 850 632 852
rect 570 843 571 845
rect 573 843 574 845
rect 570 841 574 843
rect 579 847 585 848
rect 579 845 581 847
rect 583 845 585 847
rect 579 836 585 845
rect 617 847 623 848
rect 617 845 619 847
rect 621 845 623 847
rect 617 836 623 845
rect 628 845 632 850
rect 651 854 657 855
rect 651 852 653 854
rect 655 852 657 854
rect 651 847 657 852
rect 679 855 683 858
rect 674 853 683 855
rect 694 854 695 860
rect 674 851 675 853
rect 677 851 683 853
rect 628 843 629 845
rect 631 843 632 845
rect 628 841 632 843
rect 637 845 643 846
rect 637 843 639 845
rect 641 843 643 845
rect 637 836 643 843
rect 651 845 653 847
rect 655 846 657 847
rect 674 846 678 851
rect 655 845 675 846
rect 651 844 675 845
rect 677 844 678 846
rect 651 842 678 844
rect 683 846 689 847
rect 683 844 685 846
rect 687 844 689 846
rect 683 836 689 844
rect 707 845 713 846
rect 707 843 709 845
rect 711 843 713 845
rect 707 838 713 843
rect 727 845 733 846
rect 727 843 729 845
rect 731 843 733 845
rect 707 836 709 838
rect 711 836 713 838
rect 727 838 733 843
rect 727 836 729 838
rect 731 836 733 838
rect 90 818 92 820
rect 94 818 96 820
rect 90 813 96 818
rect 110 818 112 820
rect 114 818 116 820
rect 90 811 92 813
rect 94 811 96 813
rect 90 810 96 811
rect 110 813 116 818
rect 110 811 112 813
rect 114 811 116 813
rect 110 810 116 811
rect 134 812 140 820
rect 134 810 136 812
rect 138 810 140 812
rect 134 809 140 810
rect 145 812 172 814
rect 145 810 146 812
rect 148 811 172 812
rect 148 810 168 811
rect 145 805 149 810
rect 166 809 168 810
rect 170 809 172 811
rect 180 813 186 820
rect 180 811 182 813
rect 184 811 186 813
rect 180 810 186 811
rect 191 813 195 815
rect 191 811 192 813
rect 194 811 195 813
rect 140 803 146 805
rect 148 803 149 805
rect 128 796 129 802
rect 140 801 149 803
rect 140 798 144 801
rect 166 804 172 809
rect 166 802 168 804
rect 170 802 172 804
rect 166 801 172 802
rect 191 806 195 811
rect 200 811 206 820
rect 200 809 202 811
rect 204 809 206 811
rect 200 808 206 809
rect 238 811 244 820
rect 238 809 240 811
rect 242 809 244 811
rect 238 808 244 809
rect 249 813 253 815
rect 249 811 250 813
rect 252 811 253 813
rect 191 804 192 806
rect 194 805 195 806
rect 194 804 208 805
rect 191 801 208 804
rect 132 794 144 798
rect 132 789 136 794
rect 151 793 157 794
rect 132 787 133 789
rect 135 787 136 789
rect 132 781 136 787
rect 128 775 129 781
rect 132 777 141 781
rect 204 789 208 801
rect 204 787 205 789
rect 207 787 208 789
rect 204 782 208 787
rect 196 778 208 782
rect 137 773 141 777
rect 196 774 200 778
rect 211 775 212 777
rect 180 773 200 774
rect 137 772 167 773
rect 137 770 163 772
rect 165 770 167 772
rect 180 771 182 773
rect 184 771 200 773
rect 180 770 200 771
rect 137 769 167 770
rect 249 806 253 811
rect 258 813 264 820
rect 258 811 260 813
rect 262 811 264 813
rect 258 810 264 811
rect 275 813 281 820
rect 275 811 277 813
rect 279 811 281 813
rect 275 810 281 811
rect 311 811 317 820
rect 311 809 313 811
rect 315 809 317 811
rect 311 808 317 809
rect 322 813 326 815
rect 322 811 323 813
rect 325 811 326 813
rect 249 805 250 806
rect 236 804 250 805
rect 252 804 253 806
rect 236 801 253 804
rect 236 789 240 801
rect 287 794 288 801
rect 236 787 237 789
rect 239 787 240 789
rect 236 782 240 787
rect 236 778 248 782
rect 232 775 233 777
rect 244 774 248 778
rect 273 777 277 779
rect 273 775 274 777
rect 276 775 277 777
rect 287 776 288 782
rect 244 773 264 774
rect 244 771 260 773
rect 262 771 264 773
rect 244 770 264 771
rect 108 765 114 766
rect 108 764 110 765
rect 112 764 114 765
rect 273 764 277 775
rect 322 806 326 811
rect 331 813 337 820
rect 331 811 333 813
rect 335 811 337 813
rect 331 810 337 811
rect 439 812 466 814
rect 439 811 463 812
rect 439 809 441 811
rect 443 810 463 811
rect 465 810 466 812
rect 443 809 445 810
rect 322 805 323 806
rect 309 804 323 805
rect 325 804 326 806
rect 309 801 326 804
rect 309 789 313 801
rect 439 804 445 809
rect 439 802 441 804
rect 443 802 445 804
rect 439 801 445 802
rect 462 805 466 810
rect 471 812 477 820
rect 471 810 473 812
rect 475 810 477 812
rect 471 809 477 810
rect 495 813 501 820
rect 495 811 497 813
rect 499 811 501 813
rect 495 810 501 811
rect 506 813 510 815
rect 506 811 507 813
rect 509 811 510 813
rect 462 803 463 805
rect 465 803 471 805
rect 462 801 471 803
rect 467 798 471 801
rect 467 794 479 798
rect 482 796 483 802
rect 454 793 460 794
rect 309 787 310 789
rect 312 787 313 789
rect 309 782 313 787
rect 309 778 321 782
rect 305 775 306 777
rect 317 774 321 778
rect 475 789 479 794
rect 475 787 476 789
rect 478 787 479 789
rect 475 781 479 787
rect 470 777 479 781
rect 317 773 337 774
rect 470 773 474 777
rect 482 775 483 781
rect 506 806 510 811
rect 515 811 521 820
rect 515 809 517 811
rect 519 809 521 811
rect 542 813 548 820
rect 542 811 544 813
rect 546 811 548 813
rect 542 810 548 811
rect 579 811 585 820
rect 515 808 521 809
rect 579 809 581 811
rect 583 809 585 811
rect 579 808 585 809
rect 590 813 594 815
rect 590 811 591 813
rect 593 811 594 813
rect 506 804 507 806
rect 509 805 510 806
rect 509 804 523 805
rect 506 801 523 804
rect 519 789 523 801
rect 519 787 520 789
rect 522 787 523 789
rect 519 782 523 787
rect 511 778 523 782
rect 317 771 333 773
rect 335 771 337 773
rect 317 770 337 771
rect 444 772 474 773
rect 444 770 446 772
rect 448 770 474 772
rect 444 769 474 770
rect 511 774 515 778
rect 526 775 527 777
rect 554 794 555 801
rect 495 773 515 774
rect 495 771 497 773
rect 499 771 515 773
rect 495 770 515 771
rect 540 777 544 779
rect 540 775 541 777
rect 543 775 544 777
rect 554 776 555 782
rect 540 764 544 775
rect 590 806 594 811
rect 599 813 605 820
rect 599 811 601 813
rect 603 811 605 813
rect 599 810 605 811
rect 622 813 628 820
rect 622 811 624 813
rect 626 811 628 813
rect 622 810 628 811
rect 633 813 637 815
rect 633 811 634 813
rect 636 811 637 813
rect 590 805 591 806
rect 577 804 591 805
rect 593 804 594 806
rect 577 801 594 804
rect 577 789 581 801
rect 633 806 637 811
rect 642 811 648 820
rect 642 809 644 811
rect 646 809 648 811
rect 671 813 677 820
rect 671 811 673 813
rect 675 811 677 813
rect 671 810 677 811
rect 682 813 686 815
rect 682 811 683 813
rect 685 811 686 813
rect 642 808 648 809
rect 633 804 634 806
rect 636 805 637 806
rect 636 804 650 805
rect 633 801 650 804
rect 577 787 578 789
rect 580 787 581 789
rect 577 782 581 787
rect 577 778 589 782
rect 573 775 574 777
rect 585 774 589 778
rect 646 789 650 801
rect 646 787 647 789
rect 649 787 650 789
rect 646 782 650 787
rect 638 778 650 782
rect 638 774 642 778
rect 653 775 654 777
rect 682 806 686 811
rect 691 811 697 820
rect 714 813 720 820
rect 691 809 693 811
rect 695 809 697 811
rect 691 808 697 809
rect 714 811 716 813
rect 718 811 720 813
rect 714 810 720 811
rect 725 811 731 812
rect 682 804 683 806
rect 685 805 686 806
rect 725 809 727 811
rect 729 809 731 811
rect 725 806 731 809
rect 685 804 699 805
rect 682 801 699 804
rect 695 789 699 801
rect 695 787 696 789
rect 698 787 699 789
rect 695 782 699 787
rect 687 778 699 782
rect 585 773 605 774
rect 585 771 601 773
rect 603 771 605 773
rect 585 770 605 771
rect 622 773 642 774
rect 622 771 624 773
rect 626 771 642 773
rect 622 770 642 771
rect 687 774 691 778
rect 702 775 703 777
rect 671 773 691 774
rect 671 771 673 773
rect 675 771 691 773
rect 671 770 691 771
rect 727 804 731 806
rect 729 802 731 804
rect 718 801 731 802
rect 736 811 742 820
rect 736 809 738 811
rect 740 809 742 811
rect 736 804 742 809
rect 736 802 738 804
rect 740 802 742 804
rect 736 801 742 802
rect 737 767 741 769
rect 737 765 738 767
rect 740 765 741 767
rect 737 764 741 765
rect 94 742 100 748
rect 184 743 188 748
rect 153 742 179 743
rect 94 740 96 742
rect 98 740 100 742
rect 94 739 100 740
rect 107 739 111 741
rect 107 737 108 739
rect 110 737 111 739
rect 153 740 155 742
rect 157 740 175 742
rect 177 740 179 742
rect 153 739 179 740
rect 184 741 185 743
rect 187 741 188 743
rect 184 739 188 741
rect 208 741 228 742
rect 208 739 210 741
rect 212 739 228 741
rect 81 734 85 736
rect 81 732 82 734
rect 84 732 85 734
rect 81 726 85 732
rect 107 734 111 737
rect 107 730 131 734
rect 81 722 92 726
rect 88 716 92 722
rect 127 726 131 730
rect 107 725 123 726
rect 107 723 119 725
rect 121 723 123 725
rect 107 722 123 723
rect 127 724 132 726
rect 127 722 129 724
rect 131 722 132 724
rect 107 716 111 722
rect 127 720 132 722
rect 127 718 131 720
rect 88 715 111 716
rect 88 713 90 715
rect 92 713 111 715
rect 88 712 111 713
rect 99 701 103 703
rect 99 699 100 701
rect 102 699 103 701
rect 99 694 103 699
rect 107 701 111 712
rect 115 715 131 718
rect 115 713 116 715
rect 118 714 131 715
rect 118 713 119 714
rect 115 708 119 713
rect 174 735 179 739
rect 208 738 228 739
rect 174 733 175 735
rect 177 734 200 735
rect 177 733 196 734
rect 174 732 196 733
rect 198 732 200 734
rect 174 731 200 732
rect 224 734 228 738
rect 266 742 272 748
rect 266 740 268 742
rect 270 740 272 742
rect 266 739 272 740
rect 279 739 283 741
rect 239 735 240 737
rect 224 730 236 734
rect 232 725 236 730
rect 232 723 233 725
rect 235 723 236 725
rect 115 706 116 708
rect 118 706 119 708
rect 115 704 119 706
rect 154 710 158 712
rect 154 708 155 710
rect 157 708 158 710
rect 154 703 158 708
rect 173 710 179 711
rect 173 708 175 710
rect 177 708 179 710
rect 154 701 155 703
rect 157 701 158 703
rect 107 700 140 701
rect 107 698 136 700
rect 138 698 140 700
rect 107 697 140 698
rect 99 692 100 694
rect 102 692 103 694
rect 154 692 158 701
rect 173 703 179 708
rect 232 711 236 723
rect 279 737 280 739
rect 282 737 283 739
rect 253 734 257 736
rect 253 732 254 734
rect 256 732 257 734
rect 253 726 257 732
rect 279 734 283 737
rect 279 730 303 734
rect 253 722 264 726
rect 219 708 236 711
rect 219 706 220 708
rect 222 707 236 708
rect 222 706 223 707
rect 173 701 175 703
rect 177 701 179 703
rect 173 692 179 701
rect 194 703 198 705
rect 194 701 195 703
rect 197 701 198 703
rect 194 692 198 701
rect 208 701 214 702
rect 208 699 210 701
rect 212 699 214 701
rect 208 692 214 699
rect 219 701 223 706
rect 219 699 220 701
rect 222 699 223 701
rect 219 697 223 699
rect 228 703 234 704
rect 228 701 230 703
rect 232 701 234 703
rect 228 692 234 701
rect 260 716 264 722
rect 299 726 303 730
rect 279 725 295 726
rect 279 723 291 725
rect 293 723 295 725
rect 279 722 295 723
rect 299 724 304 726
rect 299 722 301 724
rect 303 722 304 724
rect 279 716 283 722
rect 299 720 304 722
rect 299 718 303 720
rect 260 715 283 716
rect 260 713 262 715
rect 264 713 283 715
rect 260 712 283 713
rect 271 701 275 703
rect 271 699 272 701
rect 274 699 275 701
rect 271 694 275 699
rect 279 701 283 712
rect 287 715 303 718
rect 287 713 288 715
rect 290 714 303 715
rect 290 713 291 714
rect 287 708 291 713
rect 287 706 288 708
rect 290 706 291 708
rect 287 704 291 706
rect 335 737 339 748
rect 324 730 325 736
rect 335 735 336 737
rect 338 735 339 737
rect 335 733 339 735
rect 577 742 583 748
rect 535 741 555 742
rect 535 739 551 741
rect 553 739 555 741
rect 577 740 579 742
rect 581 740 583 742
rect 577 739 583 740
rect 590 739 594 741
rect 535 738 555 739
rect 324 711 325 718
rect 523 735 524 737
rect 535 734 539 738
rect 590 737 591 739
rect 593 737 594 739
rect 527 730 539 734
rect 527 725 531 730
rect 527 723 528 725
rect 530 723 531 725
rect 527 711 531 723
rect 564 734 568 736
rect 564 732 565 734
rect 567 732 568 734
rect 564 726 568 732
rect 590 734 594 737
rect 590 730 614 734
rect 564 722 575 726
rect 527 708 544 711
rect 527 707 541 708
rect 540 706 541 707
rect 543 706 544 708
rect 529 703 535 704
rect 331 701 337 702
rect 279 700 312 701
rect 279 698 308 700
rect 310 698 312 700
rect 279 697 312 698
rect 331 699 333 701
rect 335 699 337 701
rect 271 692 272 694
rect 274 692 275 694
rect 331 692 337 699
rect 529 701 531 703
rect 533 701 535 703
rect 529 692 535 701
rect 540 701 544 706
rect 571 716 575 722
rect 610 726 614 730
rect 590 725 606 726
rect 590 723 602 725
rect 604 723 606 725
rect 590 722 606 723
rect 610 724 615 726
rect 610 722 612 724
rect 614 722 615 724
rect 590 716 594 722
rect 610 720 615 722
rect 643 741 663 742
rect 643 739 645 741
rect 647 739 663 741
rect 643 738 663 739
rect 659 734 663 738
rect 674 735 675 737
rect 659 730 671 734
rect 667 725 671 730
rect 667 723 668 725
rect 670 723 671 725
rect 610 718 614 720
rect 571 715 594 716
rect 571 713 573 715
rect 575 713 594 715
rect 571 712 594 713
rect 540 699 541 701
rect 543 699 544 701
rect 540 697 544 699
rect 549 701 555 702
rect 549 699 551 701
rect 553 699 555 701
rect 549 692 555 699
rect 582 701 586 703
rect 582 699 583 701
rect 585 699 586 701
rect 582 694 586 699
rect 590 701 594 712
rect 598 715 614 718
rect 598 713 599 715
rect 601 714 614 715
rect 601 713 602 714
rect 598 708 602 713
rect 598 706 599 708
rect 601 706 602 708
rect 598 704 602 706
rect 667 711 671 723
rect 688 737 692 748
rect 688 735 689 737
rect 691 735 692 737
rect 688 733 692 735
rect 702 730 703 736
rect 716 739 720 748
rect 716 737 717 739
rect 719 737 720 739
rect 716 735 720 737
rect 654 708 671 711
rect 654 706 655 708
rect 657 707 671 708
rect 702 711 703 718
rect 657 706 658 707
rect 643 701 649 702
rect 590 700 623 701
rect 590 698 619 700
rect 621 698 623 700
rect 590 697 623 698
rect 643 699 645 701
rect 647 699 649 701
rect 582 692 583 694
rect 585 692 586 694
rect 643 692 649 699
rect 654 701 658 706
rect 654 699 655 701
rect 657 699 658 701
rect 654 697 658 699
rect 663 703 669 704
rect 663 701 665 703
rect 667 701 669 703
rect 663 692 669 701
rect 690 701 696 702
rect 690 699 692 701
rect 694 699 696 701
rect 690 692 696 699
rect 716 701 720 703
rect 716 699 717 701
rect 719 699 720 701
rect 716 694 720 699
rect 716 692 717 694
rect 719 692 720 694
rect 80 674 82 676
rect 84 674 86 676
rect 80 669 86 674
rect 80 667 82 669
rect 84 667 86 669
rect 80 666 86 667
rect 114 674 116 676
rect 118 674 120 676
rect 114 669 120 674
rect 114 667 116 669
rect 118 667 120 669
rect 114 666 120 667
rect 133 669 139 676
rect 133 667 135 669
rect 137 667 139 669
rect 133 666 139 667
rect 170 667 176 676
rect 170 665 172 667
rect 174 665 176 667
rect 170 664 176 665
rect 181 669 185 671
rect 181 667 182 669
rect 184 667 185 669
rect 181 662 185 667
rect 190 669 196 676
rect 190 667 192 669
rect 194 667 196 669
rect 190 666 196 667
rect 204 674 206 676
rect 208 674 210 676
rect 204 669 210 674
rect 204 667 206 669
rect 208 667 210 669
rect 204 666 210 667
rect 238 674 240 676
rect 242 674 244 676
rect 238 669 244 674
rect 238 667 240 669
rect 242 667 244 669
rect 238 666 244 667
rect 181 661 182 662
rect 145 650 146 657
rect 102 629 108 630
rect 102 627 104 629
rect 106 627 108 629
rect 82 622 88 623
rect 82 620 84 622
rect 86 620 88 622
rect 102 622 108 627
rect 131 633 135 635
rect 131 631 132 633
rect 134 631 135 633
rect 145 632 146 638
rect 102 620 104 622
rect 106 620 108 622
rect 131 620 135 631
rect 168 660 182 661
rect 184 660 185 662
rect 168 657 185 660
rect 168 645 172 657
rect 525 668 531 676
rect 577 674 579 676
rect 581 674 583 676
rect 525 666 527 668
rect 529 666 531 668
rect 525 665 531 666
rect 536 668 563 670
rect 536 666 537 668
rect 539 667 563 668
rect 539 666 559 667
rect 536 661 540 666
rect 557 665 559 666
rect 561 665 563 667
rect 577 669 583 674
rect 625 674 627 676
rect 629 674 631 676
rect 577 667 579 669
rect 581 667 583 669
rect 577 666 583 667
rect 602 669 606 671
rect 602 667 603 669
rect 605 667 606 669
rect 531 659 537 661
rect 539 659 540 661
rect 168 643 169 645
rect 171 643 172 645
rect 168 638 172 643
rect 168 634 180 638
rect 164 631 165 633
rect 176 630 180 634
rect 176 629 196 630
rect 176 627 192 629
rect 194 627 196 629
rect 176 626 196 627
rect 226 629 232 630
rect 226 627 228 629
rect 230 627 232 629
rect 206 622 212 623
rect 206 620 208 622
rect 210 620 212 622
rect 226 622 232 627
rect 519 652 520 658
rect 531 657 540 659
rect 531 654 535 657
rect 557 660 563 665
rect 602 662 606 667
rect 625 669 631 674
rect 625 667 627 669
rect 629 667 631 669
rect 625 666 631 667
rect 649 674 651 676
rect 653 674 655 676
rect 649 669 655 674
rect 669 674 671 676
rect 673 674 675 676
rect 649 667 651 669
rect 653 667 655 669
rect 649 666 655 667
rect 660 669 664 671
rect 660 667 661 669
rect 663 667 664 669
rect 660 663 664 667
rect 669 669 675 674
rect 720 674 721 676
rect 723 674 724 676
rect 669 667 671 669
rect 673 667 675 669
rect 683 670 716 671
rect 683 668 685 670
rect 687 668 716 670
rect 683 667 716 668
rect 669 666 675 667
rect 660 662 663 663
rect 557 658 559 660
rect 561 658 563 660
rect 557 657 563 658
rect 660 660 661 662
rect 660 658 663 660
rect 523 650 535 654
rect 523 645 527 650
rect 542 649 548 650
rect 523 643 524 645
rect 526 643 527 645
rect 523 637 527 643
rect 519 631 520 637
rect 523 633 532 637
rect 528 629 532 633
rect 651 645 652 649
rect 528 628 558 629
rect 528 626 554 628
rect 556 626 558 628
rect 528 625 558 626
rect 648 629 652 631
rect 648 627 649 629
rect 651 627 652 629
rect 226 620 228 622
rect 230 620 232 622
rect 648 622 652 627
rect 704 662 708 664
rect 704 660 705 662
rect 707 660 708 662
rect 704 655 708 660
rect 704 654 705 655
rect 692 653 705 654
rect 707 653 708 655
rect 692 650 708 653
rect 712 656 716 667
rect 720 669 724 674
rect 720 667 721 669
rect 723 667 724 669
rect 720 665 724 667
rect 712 655 735 656
rect 712 653 731 655
rect 733 653 735 655
rect 712 652 735 653
rect 692 648 696 650
rect 691 646 696 648
rect 712 646 716 652
rect 691 644 692 646
rect 694 644 696 646
rect 691 642 696 644
rect 700 645 716 646
rect 700 643 702 645
rect 704 643 716 645
rect 700 642 716 643
rect 692 638 696 642
rect 731 646 735 652
rect 731 642 742 646
rect 692 634 716 638
rect 712 631 716 634
rect 738 636 742 642
rect 738 634 739 636
rect 741 634 742 636
rect 738 632 742 634
rect 712 629 713 631
rect 715 629 716 631
rect 712 627 716 629
rect 723 628 729 629
rect 723 626 725 628
rect 727 626 729 628
rect 648 620 649 622
rect 651 620 652 622
rect 723 620 729 626
rect 94 598 100 604
rect 171 602 172 604
rect 174 602 175 604
rect 94 596 96 598
rect 98 596 100 598
rect 94 595 100 596
rect 107 595 111 597
rect 107 593 108 595
rect 110 593 111 595
rect 81 590 85 592
rect 81 588 82 590
rect 84 588 85 590
rect 81 582 85 588
rect 107 590 111 593
rect 107 586 131 590
rect 81 578 92 582
rect 88 572 92 578
rect 127 582 131 586
rect 107 581 123 582
rect 107 579 119 581
rect 121 579 123 581
rect 107 578 123 579
rect 127 580 132 582
rect 127 578 129 580
rect 131 578 132 580
rect 107 572 111 578
rect 127 576 132 578
rect 127 574 131 576
rect 88 571 111 572
rect 88 569 90 571
rect 92 569 111 571
rect 88 568 111 569
rect 99 557 103 559
rect 99 555 100 557
rect 102 555 103 557
rect 99 550 103 555
rect 107 557 111 568
rect 115 571 131 574
rect 115 569 116 571
rect 118 570 131 571
rect 118 569 119 570
rect 115 564 119 569
rect 115 562 116 564
rect 118 562 119 564
rect 115 560 119 562
rect 171 597 175 602
rect 171 595 172 597
rect 174 595 175 597
rect 171 593 175 595
rect 186 597 206 598
rect 186 595 188 597
rect 190 595 206 597
rect 186 594 206 595
rect 171 575 172 579
rect 202 590 206 594
rect 217 591 218 593
rect 202 586 214 590
rect 210 581 214 586
rect 210 579 211 581
rect 213 579 214 581
rect 160 564 163 566
rect 162 562 163 564
rect 160 561 163 562
rect 210 567 214 579
rect 197 564 214 567
rect 197 562 198 564
rect 200 563 214 564
rect 200 562 201 563
rect 148 557 154 558
rect 107 556 140 557
rect 107 554 136 556
rect 138 554 140 556
rect 107 553 140 554
rect 148 555 150 557
rect 152 555 154 557
rect 99 548 100 550
rect 102 548 103 550
rect 148 550 154 555
rect 159 557 163 561
rect 159 555 160 557
rect 162 555 163 557
rect 159 553 163 555
rect 168 557 174 558
rect 168 555 170 557
rect 172 555 174 557
rect 148 548 150 550
rect 152 548 154 550
rect 168 550 174 555
rect 168 548 170 550
rect 172 548 174 550
rect 186 557 192 558
rect 186 555 188 557
rect 190 555 192 557
rect 186 548 192 555
rect 197 557 201 562
rect 249 593 253 604
rect 238 586 239 592
rect 249 591 250 593
rect 252 591 253 593
rect 249 589 253 591
rect 520 598 524 604
rect 520 596 521 598
rect 523 596 524 598
rect 520 594 524 596
rect 562 598 566 604
rect 562 596 563 598
rect 565 596 566 598
rect 562 594 566 596
rect 592 598 622 599
rect 592 596 594 598
rect 596 596 622 598
rect 592 595 622 596
rect 238 567 239 574
rect 495 566 501 567
rect 495 564 497 566
rect 499 564 501 566
rect 197 555 198 557
rect 200 555 201 557
rect 197 553 201 555
rect 206 559 212 560
rect 206 557 208 559
rect 210 557 212 559
rect 495 559 501 564
rect 206 548 212 557
rect 245 557 251 558
rect 245 555 247 557
rect 249 555 251 557
rect 245 548 251 555
rect 495 557 497 559
rect 499 557 501 559
rect 495 548 501 557
rect 618 591 622 595
rect 562 576 563 582
rect 618 587 627 591
rect 630 587 631 593
rect 643 597 663 598
rect 643 595 645 597
rect 647 595 663 597
rect 643 594 663 595
rect 623 581 627 587
rect 623 579 624 581
rect 626 579 627 581
rect 602 574 608 575
rect 623 574 627 579
rect 615 570 627 574
rect 587 566 593 567
rect 587 564 589 566
rect 591 564 593 566
rect 587 559 593 564
rect 615 567 619 570
rect 610 565 619 567
rect 630 566 631 572
rect 659 590 663 594
rect 674 591 675 593
rect 659 586 671 590
rect 667 581 671 586
rect 667 579 668 581
rect 670 579 671 581
rect 610 563 611 565
rect 613 563 619 565
rect 587 557 589 559
rect 591 558 593 559
rect 610 558 614 563
rect 667 567 671 579
rect 688 593 692 604
rect 716 602 717 604
rect 719 602 720 604
rect 688 591 689 593
rect 691 591 692 593
rect 688 589 692 591
rect 702 586 703 592
rect 716 597 720 602
rect 716 595 717 597
rect 719 595 720 597
rect 716 593 720 595
rect 654 564 671 567
rect 654 562 655 564
rect 657 563 671 564
rect 702 567 703 574
rect 719 575 720 579
rect 657 562 658 563
rect 591 557 611 558
rect 587 556 611 557
rect 613 556 614 558
rect 587 554 614 556
rect 619 558 625 559
rect 619 556 621 558
rect 623 556 625 558
rect 619 548 625 556
rect 643 557 649 558
rect 643 555 645 557
rect 647 555 649 557
rect 643 548 649 555
rect 654 557 658 562
rect 728 564 731 566
rect 728 562 729 564
rect 728 561 731 562
rect 654 555 655 557
rect 657 555 658 557
rect 654 553 658 555
rect 663 559 669 560
rect 663 557 665 559
rect 667 557 669 559
rect 663 548 669 557
rect 690 557 696 558
rect 690 555 692 557
rect 694 555 696 557
rect 690 548 696 555
rect 717 557 723 558
rect 717 555 719 557
rect 721 555 723 557
rect 717 550 723 555
rect 728 557 732 561
rect 728 555 729 557
rect 731 555 732 557
rect 728 553 732 555
rect 737 557 743 558
rect 737 555 739 557
rect 741 555 743 557
rect 717 548 719 550
rect 721 548 723 550
rect 737 550 743 555
rect 737 548 739 550
rect 741 548 743 550
rect 80 530 82 532
rect 84 530 86 532
rect 80 525 86 530
rect 80 523 82 525
rect 84 523 86 525
rect 80 522 86 523
rect 114 530 116 532
rect 118 530 120 532
rect 114 525 120 530
rect 114 523 116 525
rect 118 523 120 525
rect 114 522 120 523
rect 131 525 137 532
rect 196 530 197 532
rect 199 530 200 532
rect 131 523 133 525
rect 135 523 137 525
rect 159 526 192 527
rect 159 524 161 526
rect 163 524 192 526
rect 159 523 192 524
rect 131 522 137 523
rect 143 506 144 513
rect 102 485 108 486
rect 102 483 104 485
rect 106 483 108 485
rect 82 478 88 479
rect 82 476 84 478
rect 86 476 88 478
rect 102 478 108 483
rect 129 489 133 491
rect 129 487 130 489
rect 132 487 133 489
rect 143 488 144 494
rect 102 476 104 478
rect 106 476 108 478
rect 129 476 133 487
rect 180 518 184 520
rect 180 516 181 518
rect 183 516 184 518
rect 180 511 184 516
rect 180 510 181 511
rect 168 509 181 510
rect 183 509 184 511
rect 168 506 184 509
rect 188 512 192 523
rect 196 525 200 530
rect 196 523 197 525
rect 199 523 200 525
rect 196 521 200 523
rect 188 511 211 512
rect 188 509 207 511
rect 209 509 211 511
rect 188 508 211 509
rect 168 504 172 506
rect 167 502 172 504
rect 188 502 192 508
rect 167 500 168 502
rect 170 500 172 502
rect 167 498 172 500
rect 176 501 192 502
rect 176 499 178 501
rect 180 499 192 501
rect 176 498 192 499
rect 168 494 172 498
rect 207 502 211 508
rect 230 523 236 532
rect 230 521 232 523
rect 234 521 236 523
rect 250 531 256 532
rect 250 529 252 531
rect 254 529 256 531
rect 250 524 256 529
rect 250 522 252 524
rect 254 522 256 524
rect 448 525 454 532
rect 500 528 504 532
rect 448 523 450 525
rect 452 523 454 525
rect 448 522 454 523
rect 250 521 256 522
rect 230 516 236 521
rect 230 514 232 516
rect 234 514 236 516
rect 230 513 236 514
rect 207 498 218 502
rect 168 490 192 494
rect 188 487 192 490
rect 214 492 218 498
rect 233 499 235 506
rect 460 506 461 513
rect 214 490 215 492
rect 217 490 218 492
rect 214 488 218 490
rect 230 488 234 490
rect 446 489 450 491
rect 188 485 189 487
rect 191 485 192 487
rect 230 486 231 488
rect 233 486 234 488
rect 446 487 447 489
rect 449 487 450 489
rect 460 488 461 494
rect 500 526 501 528
rect 503 526 504 528
rect 520 528 524 532
rect 500 524 504 526
rect 510 525 514 527
rect 510 523 511 525
rect 513 523 514 525
rect 520 526 521 528
rect 523 526 524 528
rect 572 530 573 532
rect 575 530 576 532
rect 520 524 524 526
rect 535 526 568 527
rect 535 524 537 526
rect 539 524 568 526
rect 535 523 568 524
rect 510 519 514 523
rect 493 508 498 509
rect 188 483 192 485
rect 199 484 205 485
rect 199 482 201 484
rect 203 482 205 484
rect 199 476 205 482
rect 230 476 234 486
rect 251 485 257 486
rect 251 483 253 485
rect 255 483 257 485
rect 251 476 257 483
rect 446 476 450 487
rect 493 506 494 508
rect 496 506 498 508
rect 493 505 498 506
rect 556 518 560 520
rect 556 516 557 518
rect 559 516 560 518
rect 556 511 560 516
rect 556 510 557 511
rect 544 509 557 510
rect 559 509 560 511
rect 544 506 560 509
rect 564 512 568 523
rect 572 525 576 530
rect 572 523 573 525
rect 575 523 576 525
rect 572 521 576 523
rect 603 525 609 532
rect 603 523 605 525
rect 607 523 609 525
rect 603 522 609 523
rect 614 525 618 527
rect 614 523 615 525
rect 617 523 618 525
rect 564 511 587 512
rect 564 509 583 511
rect 585 509 587 511
rect 564 508 587 509
rect 544 504 548 506
rect 543 502 548 504
rect 564 502 568 508
rect 543 500 544 502
rect 546 500 548 502
rect 543 498 548 500
rect 552 501 568 502
rect 552 499 554 501
rect 556 499 568 501
rect 552 498 568 499
rect 544 494 548 498
rect 583 502 587 508
rect 614 518 618 523
rect 623 523 629 532
rect 623 521 625 523
rect 627 521 629 523
rect 648 530 649 532
rect 651 530 652 532
rect 648 525 652 530
rect 720 530 721 532
rect 723 530 724 532
rect 683 526 716 527
rect 648 523 649 525
rect 651 523 652 525
rect 648 521 652 523
rect 683 524 685 526
rect 687 524 716 526
rect 683 523 716 524
rect 623 520 629 521
rect 614 516 615 518
rect 617 517 618 518
rect 617 516 631 517
rect 614 513 631 516
rect 583 498 594 502
rect 544 490 568 494
rect 564 487 568 490
rect 590 492 594 498
rect 590 490 591 492
rect 593 490 594 492
rect 590 488 594 490
rect 627 501 631 513
rect 627 499 628 501
rect 630 499 631 501
rect 627 494 631 499
rect 619 490 631 494
rect 564 485 565 487
rect 567 485 568 487
rect 619 486 623 490
rect 634 487 635 489
rect 603 485 623 486
rect 564 483 568 485
rect 575 484 581 485
rect 575 482 577 484
rect 579 482 581 484
rect 603 483 605 485
rect 607 483 623 485
rect 603 482 623 483
rect 575 476 581 482
rect 648 487 652 489
rect 648 485 649 487
rect 651 485 652 487
rect 648 476 652 485
rect 704 518 708 520
rect 704 516 705 518
rect 707 516 708 518
rect 704 511 708 516
rect 704 510 705 511
rect 692 509 705 510
rect 707 509 708 511
rect 692 506 708 509
rect 712 512 716 523
rect 720 525 724 530
rect 720 523 721 525
rect 723 523 724 525
rect 720 521 724 523
rect 712 511 735 512
rect 712 509 731 511
rect 733 509 735 511
rect 712 508 735 509
rect 692 504 696 506
rect 691 502 696 504
rect 712 502 716 508
rect 691 500 692 502
rect 694 500 696 502
rect 691 498 696 500
rect 700 501 716 502
rect 700 499 702 501
rect 704 499 716 501
rect 700 498 716 499
rect 692 494 696 498
rect 731 502 735 508
rect 731 498 742 502
rect 692 490 716 494
rect 712 487 716 490
rect 738 492 742 498
rect 738 490 739 492
rect 741 490 742 492
rect 738 488 742 490
rect 712 485 713 487
rect 715 485 716 487
rect 712 483 716 485
rect 723 484 729 485
rect 723 482 725 484
rect 727 482 729 484
rect 723 476 729 482
rect 18 349 24 357
rect 59 351 63 357
rect 81 355 82 357
rect 84 355 86 357
rect 81 354 86 355
rect 18 347 20 349
rect 22 347 24 349
rect 18 346 24 347
rect 48 349 55 350
rect 48 347 50 349
rect 52 347 55 349
rect 59 349 60 351
rect 62 349 63 351
rect 59 347 63 349
rect 48 346 55 347
rect 8 344 12 346
rect 8 342 9 344
rect 11 343 12 344
rect 29 344 33 346
rect 11 342 26 343
rect 8 339 26 342
rect 22 334 26 339
rect 22 332 23 334
rect 25 332 26 334
rect 22 327 26 332
rect 18 323 26 327
rect 29 342 30 344
rect 32 342 33 344
rect 18 319 22 323
rect 29 319 33 342
rect 5 318 22 319
rect 5 316 7 318
rect 9 316 22 318
rect 5 315 22 316
rect 26 318 33 319
rect 26 316 28 318
rect 30 316 33 318
rect 26 315 33 316
rect 44 334 48 336
rect 44 332 45 334
rect 47 332 48 334
rect 44 318 48 332
rect 51 325 55 346
rect 67 346 73 348
rect 67 344 70 346
rect 72 344 73 346
rect 67 342 73 344
rect 67 335 71 342
rect 58 334 71 335
rect 58 332 60 334
rect 62 332 71 334
rect 118 349 124 357
rect 159 351 163 357
rect 180 355 182 357
rect 184 355 186 357
rect 180 354 186 355
rect 92 346 97 348
rect 118 347 120 349
rect 122 347 124 349
rect 118 346 124 347
rect 148 349 155 350
rect 148 347 150 349
rect 152 347 155 349
rect 159 349 160 351
rect 162 349 163 351
rect 159 347 163 349
rect 148 346 155 347
rect 92 344 93 346
rect 95 344 97 346
rect 92 342 97 344
rect 58 331 71 332
rect 51 323 52 325
rect 54 323 55 325
rect 51 321 55 323
rect 67 327 71 331
rect 67 325 73 327
rect 67 323 70 325
rect 72 323 73 325
rect 67 321 73 323
rect 93 318 97 342
rect 108 344 112 346
rect 108 342 109 344
rect 111 343 112 344
rect 129 344 133 346
rect 111 342 126 343
rect 108 339 126 342
rect 122 334 126 339
rect 122 332 123 334
rect 125 332 126 334
rect 122 327 126 332
rect 118 323 126 327
rect 129 342 130 344
rect 132 342 133 344
rect 118 319 122 323
rect 129 319 133 342
rect 44 317 97 318
rect 44 315 93 317
rect 95 315 97 317
rect 109 315 122 319
rect 126 318 133 319
rect 126 316 128 318
rect 130 316 133 318
rect 126 315 133 316
rect 44 314 97 315
rect 144 334 148 336
rect 144 332 145 334
rect 147 332 148 334
rect 144 318 148 332
rect 151 325 155 346
rect 167 346 173 348
rect 167 344 170 346
rect 172 344 173 346
rect 167 342 173 344
rect 167 335 171 342
rect 158 334 171 335
rect 158 332 160 334
rect 162 332 171 334
rect 192 346 197 348
rect 192 344 193 346
rect 195 344 197 346
rect 192 342 197 344
rect 158 331 171 332
rect 151 323 152 325
rect 154 323 155 325
rect 151 321 155 323
rect 167 327 171 331
rect 167 325 173 327
rect 167 323 170 325
rect 172 323 173 325
rect 167 321 173 323
rect 193 318 197 342
rect 218 349 224 357
rect 259 351 263 357
rect 280 355 282 357
rect 284 355 286 357
rect 280 354 286 355
rect 218 347 220 349
rect 222 347 224 349
rect 218 346 224 347
rect 248 349 255 350
rect 248 347 250 349
rect 252 347 255 349
rect 259 349 260 351
rect 262 349 263 351
rect 259 347 263 349
rect 248 346 255 347
rect 208 344 212 346
rect 208 342 209 344
rect 211 343 212 344
rect 229 344 233 346
rect 211 342 226 343
rect 208 339 226 342
rect 222 334 226 339
rect 222 332 223 334
rect 225 332 226 334
rect 222 327 226 332
rect 218 323 226 327
rect 229 342 230 344
rect 232 342 233 344
rect 218 319 222 323
rect 229 319 233 342
rect 144 317 197 318
rect 144 315 193 317
rect 195 315 197 317
rect 205 318 222 319
rect 205 316 207 318
rect 209 316 222 318
rect 205 315 222 316
rect 226 318 233 319
rect 226 316 228 318
rect 230 316 233 318
rect 226 315 233 316
rect 144 314 197 315
rect 244 334 248 336
rect 244 332 245 334
rect 247 332 248 334
rect 244 318 248 332
rect 251 325 255 346
rect 267 346 273 348
rect 267 344 270 346
rect 272 344 273 346
rect 267 342 273 344
rect 267 335 271 342
rect 258 334 271 335
rect 258 332 260 334
rect 262 332 271 334
rect 318 349 324 357
rect 359 351 363 357
rect 380 355 382 357
rect 384 355 386 357
rect 380 354 386 355
rect 292 346 297 348
rect 318 347 320 349
rect 322 347 324 349
rect 318 346 324 347
rect 348 349 355 350
rect 348 347 350 349
rect 352 347 355 349
rect 359 349 360 351
rect 362 349 363 351
rect 359 347 363 349
rect 348 346 355 347
rect 292 344 293 346
rect 295 344 297 346
rect 292 342 297 344
rect 258 331 271 332
rect 251 323 252 325
rect 254 323 255 325
rect 251 321 255 323
rect 267 327 271 331
rect 267 325 273 327
rect 267 323 270 325
rect 272 323 273 325
rect 267 321 273 323
rect 293 318 297 342
rect 308 344 312 346
rect 308 342 309 344
rect 311 343 312 344
rect 329 344 333 346
rect 311 342 326 343
rect 308 339 326 342
rect 322 334 326 339
rect 322 332 323 334
rect 325 332 326 334
rect 322 327 326 332
rect 318 323 326 327
rect 329 342 330 344
rect 332 342 333 344
rect 318 319 322 323
rect 329 319 333 342
rect 244 317 297 318
rect 244 315 293 317
rect 295 315 297 317
rect 305 318 322 319
rect 305 316 307 318
rect 309 316 322 318
rect 305 315 322 316
rect 326 318 333 319
rect 326 316 328 318
rect 330 316 333 318
rect 326 315 333 316
rect 244 314 297 315
rect 344 334 348 336
rect 344 332 345 334
rect 347 332 348 334
rect 344 318 348 332
rect 351 325 355 346
rect 367 346 373 348
rect 418 349 424 357
rect 459 351 463 357
rect 480 355 482 357
rect 484 355 486 357
rect 480 354 486 355
rect 367 344 370 346
rect 372 344 373 346
rect 367 342 373 344
rect 367 335 371 342
rect 392 346 397 348
rect 418 347 420 349
rect 422 347 424 349
rect 418 346 424 347
rect 448 349 455 350
rect 448 347 450 349
rect 452 347 455 349
rect 459 349 460 351
rect 462 349 463 351
rect 459 347 463 349
rect 448 346 455 347
rect 392 344 393 346
rect 395 344 397 346
rect 392 342 397 344
rect 358 334 371 335
rect 358 332 360 334
rect 362 332 371 334
rect 358 331 371 332
rect 351 323 352 325
rect 354 323 355 325
rect 351 321 355 323
rect 367 327 371 331
rect 367 325 373 327
rect 367 323 370 325
rect 372 323 373 325
rect 367 321 373 323
rect 393 318 397 342
rect 408 344 412 346
rect 408 342 409 344
rect 411 343 412 344
rect 429 344 433 346
rect 411 342 426 343
rect 408 339 426 342
rect 422 334 426 339
rect 422 332 423 334
rect 425 332 426 334
rect 422 327 426 332
rect 418 323 426 327
rect 429 342 430 344
rect 432 342 433 344
rect 418 319 422 323
rect 429 319 433 342
rect 344 317 397 318
rect 344 315 393 317
rect 395 315 397 317
rect 405 318 422 319
rect 405 316 407 318
rect 409 316 422 318
rect 405 315 422 316
rect 426 318 433 319
rect 426 316 428 318
rect 430 316 433 318
rect 426 315 433 316
rect 344 314 397 315
rect 444 334 448 336
rect 444 332 445 334
rect 447 332 448 334
rect 444 318 448 332
rect 451 325 455 346
rect 467 346 473 348
rect 467 344 470 346
rect 472 344 473 346
rect 467 342 473 344
rect 467 335 471 342
rect 492 346 497 348
rect 492 344 493 346
rect 495 344 497 346
rect 492 342 497 344
rect 458 334 471 335
rect 458 332 460 334
rect 462 332 471 334
rect 458 331 471 332
rect 451 323 452 325
rect 454 323 455 325
rect 451 321 455 323
rect 467 327 471 331
rect 467 325 473 327
rect 467 323 470 325
rect 472 323 473 325
rect 467 321 473 323
rect 493 318 497 342
rect 518 349 524 357
rect 559 351 563 357
rect 580 355 582 357
rect 584 355 586 357
rect 580 354 586 355
rect 518 347 520 349
rect 522 347 524 349
rect 518 346 524 347
rect 548 349 555 350
rect 548 347 550 349
rect 552 347 555 349
rect 559 349 560 351
rect 562 349 563 351
rect 559 347 563 349
rect 548 346 555 347
rect 508 344 512 346
rect 508 342 509 344
rect 511 343 512 344
rect 529 344 533 346
rect 511 342 526 343
rect 508 339 526 342
rect 522 334 526 339
rect 522 332 523 334
rect 525 332 526 334
rect 522 327 526 332
rect 518 323 526 327
rect 529 342 530 344
rect 532 342 533 344
rect 518 319 522 323
rect 529 319 533 342
rect 444 317 497 318
rect 444 315 493 317
rect 495 315 497 317
rect 505 318 522 319
rect 505 316 507 318
rect 509 316 522 318
rect 505 315 522 316
rect 526 318 533 319
rect 526 316 528 318
rect 530 316 533 318
rect 526 315 533 316
rect 444 314 497 315
rect 544 334 548 336
rect 544 332 545 334
rect 547 332 548 334
rect 544 318 548 332
rect 551 325 555 346
rect 567 346 573 348
rect 567 344 570 346
rect 572 344 573 346
rect 567 342 573 344
rect 567 335 571 342
rect 592 346 597 348
rect 592 344 593 346
rect 595 344 597 346
rect 592 342 597 344
rect 558 334 571 335
rect 558 332 560 334
rect 562 332 571 334
rect 558 331 571 332
rect 551 323 552 325
rect 554 323 555 325
rect 551 321 555 323
rect 567 327 571 331
rect 567 325 573 327
rect 567 323 570 325
rect 572 323 573 325
rect 567 321 573 323
rect 593 318 597 342
rect 618 349 624 357
rect 659 351 663 357
rect 680 355 682 357
rect 684 355 686 357
rect 680 354 686 355
rect 618 347 620 349
rect 622 347 624 349
rect 618 346 624 347
rect 648 349 655 350
rect 648 347 650 349
rect 652 347 655 349
rect 659 349 660 351
rect 662 349 663 351
rect 659 347 663 349
rect 648 346 655 347
rect 608 344 612 346
rect 608 342 609 344
rect 611 343 612 344
rect 629 344 633 346
rect 611 342 626 343
rect 608 339 626 342
rect 622 334 626 339
rect 622 332 623 334
rect 625 332 626 334
rect 622 327 626 332
rect 618 323 626 327
rect 629 342 630 344
rect 632 342 633 344
rect 618 319 622 323
rect 629 319 633 342
rect 544 317 597 318
rect 544 315 593 317
rect 595 315 597 317
rect 605 318 622 319
rect 605 316 607 318
rect 609 316 622 318
rect 605 315 622 316
rect 626 318 633 319
rect 626 316 628 318
rect 630 316 633 318
rect 626 315 633 316
rect 544 314 597 315
rect 644 334 648 336
rect 644 332 645 334
rect 647 332 648 334
rect 644 318 648 332
rect 651 325 655 346
rect 667 346 673 348
rect 667 344 670 346
rect 672 344 673 346
rect 667 342 673 344
rect 667 335 671 342
rect 692 346 697 348
rect 692 344 693 346
rect 695 344 697 346
rect 692 342 697 344
rect 658 334 671 335
rect 658 332 660 334
rect 662 332 671 334
rect 658 331 671 332
rect 651 323 652 325
rect 654 323 655 325
rect 651 321 655 323
rect 667 327 671 331
rect 667 325 673 327
rect 667 323 670 325
rect 672 323 673 325
rect 667 321 673 323
rect 693 318 697 342
rect 718 349 724 357
rect 759 351 763 357
rect 780 355 782 357
rect 784 355 786 357
rect 780 354 786 355
rect 718 347 720 349
rect 722 347 724 349
rect 718 346 724 347
rect 748 349 755 350
rect 748 347 750 349
rect 752 347 755 349
rect 759 349 760 351
rect 762 349 763 351
rect 759 347 763 349
rect 748 346 755 347
rect 708 344 712 346
rect 708 342 709 344
rect 711 343 712 344
rect 729 344 733 346
rect 711 342 726 343
rect 708 339 726 342
rect 722 334 726 339
rect 722 332 723 334
rect 725 332 726 334
rect 722 327 726 332
rect 718 323 726 327
rect 729 342 730 344
rect 732 342 733 344
rect 718 319 722 323
rect 729 319 733 342
rect 644 317 697 318
rect 644 315 693 317
rect 695 315 697 317
rect 705 318 722 319
rect 705 316 707 318
rect 709 316 722 318
rect 705 315 722 316
rect 726 318 733 319
rect 726 316 728 318
rect 730 316 733 318
rect 726 315 733 316
rect 644 314 697 315
rect 744 334 748 336
rect 744 332 745 334
rect 747 332 748 334
rect 744 318 748 332
rect 751 325 755 346
rect 767 346 773 348
rect 767 344 770 346
rect 772 344 773 346
rect 767 342 773 344
rect 767 335 771 342
rect 792 346 797 348
rect 792 344 793 346
rect 795 344 797 346
rect 792 342 797 344
rect 758 334 771 335
rect 758 332 760 334
rect 762 332 771 334
rect 758 331 771 332
rect 751 323 752 325
rect 754 323 755 325
rect 751 321 755 323
rect 767 327 771 331
rect 767 325 773 327
rect 767 323 770 325
rect 772 323 773 325
rect 767 321 773 323
rect 793 318 797 342
rect 744 317 797 318
rect 744 315 793 317
rect 795 315 797 317
rect 744 314 797 315
rect 16 310 22 311
rect 16 308 18 310
rect 20 308 22 310
rect 16 301 22 308
rect 116 310 122 311
rect 60 309 66 310
rect 60 307 62 309
rect 64 307 66 309
rect 60 301 66 307
rect 79 309 85 310
rect 79 307 81 309
rect 83 307 85 309
rect 79 301 85 307
rect 116 308 118 310
rect 120 308 122 310
rect 116 301 122 308
rect 216 310 222 311
rect 160 309 166 310
rect 160 307 162 309
rect 164 307 166 309
rect 160 301 166 307
rect 179 309 185 310
rect 179 307 181 309
rect 183 307 185 309
rect 179 301 185 307
rect 216 308 218 310
rect 220 308 222 310
rect 216 301 222 308
rect 316 310 322 311
rect 260 309 266 310
rect 260 307 262 309
rect 264 307 266 309
rect 260 301 266 307
rect 279 309 285 310
rect 279 307 281 309
rect 283 307 285 309
rect 279 301 285 307
rect 316 308 318 310
rect 320 308 322 310
rect 316 301 322 308
rect 416 310 422 311
rect 360 309 366 310
rect 360 307 362 309
rect 364 307 366 309
rect 360 301 366 307
rect 379 309 385 310
rect 379 307 381 309
rect 383 307 385 309
rect 379 301 385 307
rect 416 308 418 310
rect 420 308 422 310
rect 416 301 422 308
rect 516 310 522 311
rect 460 309 466 310
rect 460 307 462 309
rect 464 307 466 309
rect 460 301 466 307
rect 479 309 485 310
rect 479 307 481 309
rect 483 307 485 309
rect 479 301 485 307
rect 516 308 518 310
rect 520 308 522 310
rect 516 301 522 308
rect 616 310 622 311
rect 560 309 566 310
rect 560 307 562 309
rect 564 307 566 309
rect 560 301 566 307
rect 579 309 585 310
rect 579 307 581 309
rect 583 307 585 309
rect 579 301 585 307
rect 616 308 618 310
rect 620 308 622 310
rect 616 301 622 308
rect 716 310 722 311
rect 660 309 666 310
rect 660 307 662 309
rect 664 307 666 309
rect 660 301 666 307
rect 679 309 685 310
rect 679 307 681 309
rect 683 307 685 309
rect 679 301 685 307
rect 716 308 718 310
rect 720 308 722 310
rect 716 301 722 308
rect 760 309 766 310
rect 760 307 762 309
rect 764 307 766 309
rect 760 301 766 307
rect 779 309 785 310
rect 779 307 781 309
rect 783 307 785 309
rect 779 301 785 307
rect 17 279 23 285
rect 17 277 19 279
rect 21 277 23 279
rect 17 276 23 277
rect 36 279 42 285
rect 36 277 38 279
rect 40 277 42 279
rect 36 276 42 277
rect 80 278 86 285
rect 80 276 82 278
rect 84 276 86 278
rect 117 279 123 285
rect 117 277 119 279
rect 121 277 123 279
rect 117 276 123 277
rect 136 279 142 285
rect 136 277 138 279
rect 140 277 142 279
rect 136 276 142 277
rect 80 275 86 276
rect 180 278 186 285
rect 180 276 182 278
rect 184 276 186 278
rect 217 279 223 285
rect 217 277 219 279
rect 221 277 223 279
rect 217 276 223 277
rect 236 279 242 285
rect 236 277 238 279
rect 240 277 242 279
rect 236 276 242 277
rect 180 275 186 276
rect 280 278 286 285
rect 280 276 282 278
rect 284 276 286 278
rect 317 279 323 285
rect 317 277 319 279
rect 321 277 323 279
rect 317 276 323 277
rect 336 279 342 285
rect 336 277 338 279
rect 340 277 342 279
rect 336 276 342 277
rect 280 275 286 276
rect 380 278 386 285
rect 380 276 382 278
rect 384 276 386 278
rect 419 279 425 285
rect 419 277 421 279
rect 423 277 425 279
rect 419 276 425 277
rect 438 279 444 285
rect 438 277 440 279
rect 442 277 444 279
rect 438 276 444 277
rect 380 275 386 276
rect 482 278 488 285
rect 482 276 484 278
rect 486 276 488 278
rect 519 279 525 285
rect 519 277 521 279
rect 523 277 525 279
rect 519 276 525 277
rect 538 279 544 285
rect 538 277 540 279
rect 542 277 544 279
rect 538 276 544 277
rect 482 275 488 276
rect 582 278 588 285
rect 582 276 584 278
rect 586 276 588 278
rect 619 279 625 285
rect 619 277 621 279
rect 623 277 625 279
rect 619 276 625 277
rect 638 279 644 285
rect 638 277 640 279
rect 642 277 644 279
rect 638 276 644 277
rect 582 275 588 276
rect 682 278 688 285
rect 682 276 684 278
rect 686 276 688 278
rect 719 279 725 285
rect 719 277 721 279
rect 723 277 725 279
rect 719 276 725 277
rect 738 279 744 285
rect 738 277 740 279
rect 742 277 744 279
rect 738 276 744 277
rect 682 275 688 276
rect 782 278 788 285
rect 782 276 784 278
rect 786 276 788 278
rect 782 275 788 276
rect 5 271 58 272
rect 5 269 7 271
rect 9 269 58 271
rect 5 268 58 269
rect 5 244 9 268
rect 29 263 35 265
rect 29 261 30 263
rect 32 261 35 263
rect 29 259 35 261
rect 31 255 35 259
rect 47 263 51 265
rect 47 261 48 263
rect 50 261 51 263
rect 31 254 44 255
rect 31 252 40 254
rect 42 252 44 254
rect 31 251 44 252
rect 5 242 10 244
rect 5 240 7 242
rect 9 240 10 242
rect 5 238 10 240
rect 31 244 35 251
rect 29 242 35 244
rect 29 240 30 242
rect 32 240 35 242
rect 29 238 35 240
rect 47 240 51 261
rect 54 254 58 268
rect 54 252 55 254
rect 57 252 58 254
rect 54 250 58 252
rect 105 271 158 272
rect 69 270 76 271
rect 69 268 72 270
rect 74 268 76 270
rect 69 267 76 268
rect 80 270 96 271
rect 80 268 93 270
rect 95 268 96 270
rect 80 267 96 268
rect 105 269 107 271
rect 109 269 158 271
rect 105 268 158 269
rect 69 244 73 267
rect 80 263 84 267
rect 69 242 70 244
rect 72 242 73 244
rect 76 259 84 263
rect 76 254 80 259
rect 76 252 77 254
rect 79 252 80 254
rect 76 247 80 252
rect 76 244 94 247
rect 76 243 91 244
rect 69 240 73 242
rect 90 242 91 243
rect 93 242 94 244
rect 90 240 94 242
rect 47 239 54 240
rect 39 237 43 239
rect 39 235 40 237
rect 42 235 43 237
rect 47 237 50 239
rect 52 237 54 239
rect 47 236 54 237
rect 78 239 84 240
rect 78 237 80 239
rect 82 237 84 239
rect 16 231 22 232
rect 16 229 18 231
rect 20 229 22 231
rect 39 229 43 235
rect 78 229 84 237
rect 105 244 109 268
rect 129 263 135 265
rect 129 261 130 263
rect 132 261 135 263
rect 129 259 135 261
rect 131 255 135 259
rect 147 263 151 265
rect 147 261 148 263
rect 150 261 151 263
rect 131 254 144 255
rect 131 252 140 254
rect 142 252 144 254
rect 131 251 144 252
rect 105 242 110 244
rect 105 240 107 242
rect 109 240 110 242
rect 105 238 110 240
rect 131 244 135 251
rect 129 242 135 244
rect 129 240 130 242
rect 132 240 135 242
rect 129 238 135 240
rect 147 240 151 261
rect 154 254 158 268
rect 154 252 155 254
rect 157 252 158 254
rect 154 250 158 252
rect 205 271 258 272
rect 169 270 176 271
rect 169 268 172 270
rect 174 268 176 270
rect 169 267 176 268
rect 180 270 197 271
rect 180 268 193 270
rect 195 268 197 270
rect 180 267 197 268
rect 205 269 207 271
rect 209 269 258 271
rect 205 268 258 269
rect 169 244 173 267
rect 180 263 184 267
rect 169 242 170 244
rect 172 242 173 244
rect 176 259 184 263
rect 176 254 180 259
rect 176 252 177 254
rect 179 252 180 254
rect 176 247 180 252
rect 176 244 194 247
rect 176 243 191 244
rect 169 240 173 242
rect 190 242 191 243
rect 193 242 194 244
rect 190 240 194 242
rect 205 244 209 268
rect 229 263 235 265
rect 229 261 230 263
rect 232 261 235 263
rect 229 259 235 261
rect 231 255 235 259
rect 247 263 251 265
rect 247 261 248 263
rect 250 261 251 263
rect 231 254 244 255
rect 231 252 240 254
rect 242 252 244 254
rect 231 251 244 252
rect 205 242 210 244
rect 205 240 207 242
rect 209 240 210 242
rect 147 239 154 240
rect 139 237 143 239
rect 139 235 140 237
rect 142 235 143 237
rect 147 237 150 239
rect 152 237 154 239
rect 147 236 154 237
rect 178 239 184 240
rect 178 237 180 239
rect 182 237 184 239
rect 205 238 210 240
rect 231 244 235 251
rect 229 242 235 244
rect 229 240 230 242
rect 232 240 235 242
rect 116 231 122 232
rect 116 229 118 231
rect 120 229 122 231
rect 139 229 143 235
rect 178 229 184 237
rect 229 238 235 240
rect 247 240 251 261
rect 254 254 258 268
rect 254 252 255 254
rect 257 252 258 254
rect 254 250 258 252
rect 280 271 297 272
rect 269 270 276 271
rect 269 268 272 270
rect 274 268 276 270
rect 269 267 276 268
rect 280 269 293 271
rect 295 269 297 271
rect 280 268 297 269
rect 305 271 358 272
rect 305 269 307 271
rect 309 269 358 271
rect 305 268 358 269
rect 269 244 273 267
rect 280 263 284 268
rect 269 242 270 244
rect 272 242 273 244
rect 276 259 284 263
rect 276 254 280 259
rect 276 252 277 254
rect 279 252 280 254
rect 276 247 280 252
rect 276 244 294 247
rect 276 243 291 244
rect 269 240 273 242
rect 290 242 291 243
rect 293 242 294 244
rect 290 240 294 242
rect 305 244 309 268
rect 329 263 335 265
rect 329 261 330 263
rect 332 261 335 263
rect 329 259 335 261
rect 331 255 335 259
rect 347 263 351 265
rect 347 261 348 263
rect 350 261 351 263
rect 331 254 344 255
rect 331 252 340 254
rect 342 252 344 254
rect 331 251 344 252
rect 305 242 310 244
rect 305 240 307 242
rect 309 240 310 242
rect 247 239 254 240
rect 239 237 243 239
rect 239 235 240 237
rect 242 235 243 237
rect 247 237 250 239
rect 252 237 254 239
rect 247 236 254 237
rect 278 239 284 240
rect 278 237 280 239
rect 282 237 284 239
rect 305 238 310 240
rect 331 244 335 251
rect 329 242 335 244
rect 329 240 330 242
rect 332 240 335 242
rect 216 231 222 232
rect 216 229 218 231
rect 220 229 222 231
rect 239 229 243 235
rect 278 229 284 237
rect 329 238 335 240
rect 347 240 351 261
rect 354 254 358 268
rect 354 252 355 254
rect 357 252 358 254
rect 354 250 358 252
rect 407 271 460 272
rect 369 270 376 271
rect 369 268 372 270
rect 374 268 376 270
rect 369 267 376 268
rect 380 270 397 271
rect 380 268 393 270
rect 395 268 397 270
rect 380 267 397 268
rect 407 269 409 271
rect 411 269 460 271
rect 407 268 460 269
rect 369 244 373 267
rect 380 263 384 267
rect 369 242 370 244
rect 372 242 373 244
rect 376 259 384 263
rect 376 254 380 259
rect 376 252 377 254
rect 379 252 380 254
rect 376 247 380 252
rect 376 244 394 247
rect 376 243 391 244
rect 369 240 373 242
rect 390 242 391 243
rect 393 242 394 244
rect 390 240 394 242
rect 347 239 354 240
rect 339 237 343 239
rect 339 235 340 237
rect 342 235 343 237
rect 347 237 350 239
rect 352 237 354 239
rect 347 236 354 237
rect 378 239 384 240
rect 378 237 380 239
rect 382 237 384 239
rect 316 231 322 232
rect 316 229 318 231
rect 320 229 322 231
rect 339 229 343 235
rect 378 229 384 237
rect 407 244 411 268
rect 431 263 437 265
rect 431 261 432 263
rect 434 261 437 263
rect 431 259 437 261
rect 433 255 437 259
rect 449 263 453 265
rect 449 261 450 263
rect 452 261 453 263
rect 433 254 446 255
rect 433 252 442 254
rect 444 252 446 254
rect 433 251 446 252
rect 407 242 412 244
rect 407 240 409 242
rect 411 240 412 242
rect 407 238 412 240
rect 433 244 437 251
rect 431 242 437 244
rect 431 240 432 242
rect 434 240 437 242
rect 431 238 437 240
rect 449 240 453 261
rect 456 254 460 268
rect 456 252 457 254
rect 459 252 460 254
rect 456 250 460 252
rect 482 271 499 272
rect 471 270 478 271
rect 471 268 474 270
rect 476 268 478 270
rect 471 267 478 268
rect 482 269 495 271
rect 497 269 499 271
rect 482 268 499 269
rect 507 271 560 272
rect 507 269 509 271
rect 511 269 560 271
rect 507 268 560 269
rect 471 244 475 267
rect 482 263 486 268
rect 471 242 472 244
rect 474 242 475 244
rect 478 259 486 263
rect 478 254 482 259
rect 478 252 479 254
rect 481 252 482 254
rect 478 247 482 252
rect 478 244 496 247
rect 478 243 493 244
rect 471 240 475 242
rect 492 242 493 243
rect 495 242 496 244
rect 492 240 496 242
rect 507 244 511 268
rect 531 263 537 265
rect 531 261 532 263
rect 534 261 537 263
rect 531 259 537 261
rect 533 255 537 259
rect 549 263 553 265
rect 549 261 550 263
rect 552 261 553 263
rect 533 254 546 255
rect 533 252 542 254
rect 544 252 546 254
rect 533 251 546 252
rect 507 242 512 244
rect 507 240 509 242
rect 511 240 512 242
rect 449 239 456 240
rect 441 237 445 239
rect 441 235 442 237
rect 444 235 445 237
rect 449 237 452 239
rect 454 237 456 239
rect 449 236 456 237
rect 480 239 486 240
rect 480 237 482 239
rect 484 237 486 239
rect 507 238 512 240
rect 533 244 537 251
rect 531 242 537 244
rect 531 240 532 242
rect 534 240 537 242
rect 418 231 424 232
rect 418 229 420 231
rect 422 229 424 231
rect 441 229 445 235
rect 480 229 486 237
rect 531 238 537 240
rect 549 240 553 261
rect 556 254 560 268
rect 556 252 557 254
rect 559 252 560 254
rect 556 250 560 252
rect 607 271 660 272
rect 571 270 578 271
rect 571 268 574 270
rect 576 268 578 270
rect 571 267 578 268
rect 582 270 599 271
rect 582 268 595 270
rect 597 268 599 270
rect 582 267 599 268
rect 607 269 609 271
rect 611 269 660 271
rect 607 268 660 269
rect 571 244 575 267
rect 582 263 586 267
rect 571 242 572 244
rect 574 242 575 244
rect 578 259 586 263
rect 578 254 582 259
rect 578 252 579 254
rect 581 252 582 254
rect 578 247 582 252
rect 578 244 596 247
rect 578 243 593 244
rect 571 240 575 242
rect 592 242 593 243
rect 595 242 596 244
rect 592 240 596 242
rect 607 244 611 268
rect 631 263 637 265
rect 631 261 632 263
rect 634 261 637 263
rect 631 259 637 261
rect 633 255 637 259
rect 649 263 653 265
rect 649 261 650 263
rect 652 261 653 263
rect 633 254 646 255
rect 633 252 642 254
rect 644 252 646 254
rect 633 251 646 252
rect 607 242 612 244
rect 607 240 609 242
rect 611 240 612 242
rect 549 239 556 240
rect 541 237 545 239
rect 541 235 542 237
rect 544 235 545 237
rect 549 237 552 239
rect 554 237 556 239
rect 549 236 556 237
rect 580 239 586 240
rect 580 237 582 239
rect 584 237 586 239
rect 607 238 612 240
rect 633 244 637 251
rect 631 242 637 244
rect 631 240 632 242
rect 634 240 637 242
rect 518 231 524 232
rect 518 229 520 231
rect 522 229 524 231
rect 541 229 545 235
rect 580 229 586 237
rect 631 238 637 240
rect 649 240 653 261
rect 656 254 660 268
rect 656 252 657 254
rect 659 252 660 254
rect 656 250 660 252
rect 682 271 699 272
rect 671 270 678 271
rect 671 268 674 270
rect 676 268 678 270
rect 671 267 678 268
rect 682 269 695 271
rect 697 269 699 271
rect 682 268 699 269
rect 707 271 760 272
rect 707 269 709 271
rect 711 269 760 271
rect 707 268 760 269
rect 671 244 675 267
rect 682 263 686 268
rect 671 242 672 244
rect 674 242 675 244
rect 678 259 686 263
rect 678 254 682 259
rect 678 252 679 254
rect 681 252 682 254
rect 678 247 682 252
rect 678 244 696 247
rect 678 243 693 244
rect 671 240 675 242
rect 692 242 693 243
rect 695 242 696 244
rect 692 240 696 242
rect 707 244 711 268
rect 731 263 737 265
rect 731 261 732 263
rect 734 261 737 263
rect 731 259 737 261
rect 733 255 737 259
rect 749 263 753 265
rect 749 261 750 263
rect 752 261 753 263
rect 733 254 746 255
rect 733 252 742 254
rect 744 252 746 254
rect 733 251 746 252
rect 707 242 712 244
rect 707 240 709 242
rect 711 240 712 242
rect 649 239 656 240
rect 641 237 645 239
rect 641 235 642 237
rect 644 235 645 237
rect 649 237 652 239
rect 654 237 656 239
rect 649 236 656 237
rect 680 239 686 240
rect 680 237 682 239
rect 684 237 686 239
rect 707 238 712 240
rect 733 244 737 251
rect 731 242 737 244
rect 731 240 732 242
rect 734 240 737 242
rect 618 231 624 232
rect 618 229 620 231
rect 622 229 624 231
rect 641 229 645 235
rect 680 229 686 237
rect 731 238 737 240
rect 749 240 753 261
rect 756 254 760 268
rect 756 252 757 254
rect 759 252 760 254
rect 756 250 760 252
rect 771 270 778 271
rect 771 268 774 270
rect 776 268 778 270
rect 771 267 778 268
rect 782 270 799 271
rect 782 268 795 270
rect 797 268 799 270
rect 782 267 799 268
rect 771 244 775 267
rect 782 263 786 267
rect 771 242 772 244
rect 774 242 775 244
rect 778 259 786 263
rect 778 254 782 259
rect 778 252 779 254
rect 781 252 782 254
rect 778 247 782 252
rect 778 244 796 247
rect 778 243 793 244
rect 771 240 775 242
rect 792 242 793 243
rect 795 242 796 244
rect 792 240 796 242
rect 749 239 756 240
rect 741 237 745 239
rect 741 235 742 237
rect 744 235 745 237
rect 749 237 752 239
rect 754 237 756 239
rect 749 236 756 237
rect 780 239 786 240
rect 780 237 782 239
rect 784 237 786 239
rect 718 231 724 232
rect 718 229 720 231
rect 722 229 724 231
rect 741 229 745 235
rect 780 229 786 237
rect 16 211 18 213
rect 20 211 22 213
rect 16 210 22 211
rect 39 207 43 213
rect 5 202 10 204
rect 5 200 7 202
rect 9 200 10 202
rect 5 198 10 200
rect 39 205 40 207
rect 42 205 43 207
rect 5 174 9 198
rect 29 202 35 204
rect 39 203 43 205
rect 47 205 54 206
rect 47 203 50 205
rect 52 203 54 205
rect 29 200 30 202
rect 32 200 35 202
rect 29 198 35 200
rect 31 191 35 198
rect 47 202 54 203
rect 78 205 84 213
rect 116 211 118 213
rect 120 211 122 213
rect 116 210 122 211
rect 139 207 143 213
rect 78 203 80 205
rect 82 203 84 205
rect 78 202 84 203
rect 31 190 44 191
rect 31 188 40 190
rect 42 188 44 190
rect 31 187 44 188
rect 31 183 35 187
rect 29 181 35 183
rect 29 179 30 181
rect 32 179 35 181
rect 29 177 35 179
rect 47 181 51 202
rect 47 179 48 181
rect 50 179 51 181
rect 47 177 51 179
rect 54 190 58 192
rect 54 188 55 190
rect 57 188 58 190
rect 54 174 58 188
rect 5 173 58 174
rect 5 171 7 173
rect 9 171 58 173
rect 5 170 58 171
rect 69 200 73 202
rect 69 198 70 200
rect 72 198 73 200
rect 90 200 94 202
rect 90 199 91 200
rect 69 175 73 198
rect 76 198 91 199
rect 93 198 94 200
rect 76 195 94 198
rect 76 190 80 195
rect 76 188 77 190
rect 79 188 80 190
rect 76 183 80 188
rect 105 202 110 204
rect 105 200 107 202
rect 109 200 110 202
rect 105 198 110 200
rect 139 205 140 207
rect 142 205 143 207
rect 76 179 84 183
rect 80 175 84 179
rect 69 174 76 175
rect 69 172 72 174
rect 74 172 76 174
rect 69 171 76 172
rect 80 174 97 175
rect 80 172 93 174
rect 95 172 97 174
rect 80 171 97 172
rect 105 174 109 198
rect 129 202 135 204
rect 139 203 143 205
rect 147 205 154 206
rect 147 203 150 205
rect 152 203 154 205
rect 129 200 130 202
rect 132 200 135 202
rect 129 198 135 200
rect 131 191 135 198
rect 147 202 154 203
rect 178 205 184 213
rect 216 211 218 213
rect 220 211 222 213
rect 216 210 222 211
rect 239 207 243 213
rect 178 203 180 205
rect 182 203 184 205
rect 178 202 184 203
rect 205 202 210 204
rect 131 190 144 191
rect 131 188 140 190
rect 142 188 144 190
rect 131 187 144 188
rect 131 183 135 187
rect 129 181 135 183
rect 129 179 130 181
rect 132 179 135 181
rect 129 177 135 179
rect 147 181 151 202
rect 147 179 148 181
rect 150 179 151 181
rect 147 177 151 179
rect 154 190 158 192
rect 154 188 155 190
rect 157 188 158 190
rect 154 174 158 188
rect 105 173 158 174
rect 105 171 107 173
rect 109 171 158 173
rect 105 170 158 171
rect 169 200 173 202
rect 169 198 170 200
rect 172 198 173 200
rect 190 200 194 202
rect 190 199 191 200
rect 169 175 173 198
rect 176 198 191 199
rect 193 198 194 200
rect 176 195 194 198
rect 205 200 207 202
rect 209 200 210 202
rect 205 198 210 200
rect 239 205 240 207
rect 242 205 243 207
rect 176 190 180 195
rect 176 188 177 190
rect 179 188 180 190
rect 176 183 180 188
rect 176 179 184 183
rect 180 175 184 179
rect 169 174 176 175
rect 169 172 172 174
rect 174 172 176 174
rect 169 171 176 172
rect 180 174 197 175
rect 180 172 193 174
rect 195 172 197 174
rect 180 171 197 172
rect 205 174 209 198
rect 229 202 235 204
rect 239 203 243 205
rect 247 205 254 206
rect 247 203 250 205
rect 252 203 254 205
rect 229 200 230 202
rect 232 200 235 202
rect 229 198 235 200
rect 231 191 235 198
rect 247 202 254 203
rect 278 205 284 213
rect 316 211 318 213
rect 320 211 322 213
rect 316 210 322 211
rect 339 207 343 213
rect 278 203 280 205
rect 282 203 284 205
rect 278 202 284 203
rect 231 190 244 191
rect 231 188 240 190
rect 242 188 244 190
rect 231 187 244 188
rect 231 183 235 187
rect 229 181 235 183
rect 229 179 230 181
rect 232 179 235 181
rect 229 177 235 179
rect 247 181 251 202
rect 247 179 248 181
rect 250 179 251 181
rect 247 177 251 179
rect 254 190 258 192
rect 254 188 255 190
rect 257 188 258 190
rect 254 174 258 188
rect 205 173 258 174
rect 205 171 207 173
rect 209 171 258 173
rect 205 170 258 171
rect 269 200 273 202
rect 269 198 270 200
rect 272 198 273 200
rect 290 200 294 202
rect 290 199 291 200
rect 269 175 273 198
rect 276 198 291 199
rect 293 198 294 200
rect 276 195 294 198
rect 276 190 280 195
rect 276 188 277 190
rect 279 188 280 190
rect 276 183 280 188
rect 305 202 310 204
rect 305 200 307 202
rect 309 200 310 202
rect 305 198 310 200
rect 339 205 340 207
rect 342 205 343 207
rect 276 179 284 183
rect 280 175 284 179
rect 269 174 276 175
rect 269 172 272 174
rect 274 172 276 174
rect 269 171 276 172
rect 280 174 297 175
rect 280 172 293 174
rect 295 172 297 174
rect 280 171 297 172
rect 305 174 309 198
rect 329 202 335 204
rect 339 203 343 205
rect 347 205 354 206
rect 347 203 350 205
rect 352 203 354 205
rect 329 200 330 202
rect 332 200 335 202
rect 329 198 335 200
rect 331 191 335 198
rect 347 202 354 203
rect 378 205 384 213
rect 418 211 420 213
rect 422 211 424 213
rect 418 210 424 211
rect 441 207 445 213
rect 378 203 380 205
rect 382 203 384 205
rect 378 202 384 203
rect 331 190 344 191
rect 331 188 340 190
rect 342 188 344 190
rect 331 187 344 188
rect 331 183 335 187
rect 329 181 335 183
rect 329 179 330 181
rect 332 179 335 181
rect 329 177 335 179
rect 347 181 351 202
rect 347 179 348 181
rect 350 179 351 181
rect 347 177 351 179
rect 354 190 358 192
rect 354 188 355 190
rect 357 188 358 190
rect 354 174 358 188
rect 305 173 358 174
rect 305 171 307 173
rect 309 171 358 173
rect 305 170 358 171
rect 369 200 373 202
rect 369 198 370 200
rect 372 198 373 200
rect 390 200 394 202
rect 390 199 391 200
rect 369 175 373 198
rect 376 198 391 199
rect 393 198 394 200
rect 376 195 394 198
rect 376 190 380 195
rect 376 188 377 190
rect 379 188 380 190
rect 376 183 380 188
rect 407 202 412 204
rect 407 200 409 202
rect 411 200 412 202
rect 407 198 412 200
rect 441 205 442 207
rect 444 205 445 207
rect 376 179 384 183
rect 380 175 384 179
rect 369 174 376 175
rect 369 172 372 174
rect 374 172 376 174
rect 369 171 376 172
rect 380 174 397 175
rect 380 172 393 174
rect 395 172 397 174
rect 380 171 397 172
rect 407 174 411 198
rect 431 202 437 204
rect 441 203 445 205
rect 449 205 456 206
rect 449 203 452 205
rect 454 203 456 205
rect 431 200 432 202
rect 434 200 437 202
rect 431 198 437 200
rect 433 191 437 198
rect 449 202 456 203
rect 480 205 486 213
rect 518 211 520 213
rect 522 211 524 213
rect 518 210 524 211
rect 541 207 545 213
rect 480 203 482 205
rect 484 203 486 205
rect 480 202 486 203
rect 507 202 512 204
rect 433 190 446 191
rect 433 188 442 190
rect 444 188 446 190
rect 433 187 446 188
rect 433 183 437 187
rect 431 181 437 183
rect 431 179 432 181
rect 434 179 437 181
rect 431 177 437 179
rect 449 181 453 202
rect 449 179 450 181
rect 452 179 453 181
rect 449 177 453 179
rect 456 190 460 192
rect 456 188 457 190
rect 459 188 460 190
rect 456 174 460 188
rect 407 173 460 174
rect 407 171 409 173
rect 411 171 460 173
rect 407 170 460 171
rect 471 200 475 202
rect 471 198 472 200
rect 474 198 475 200
rect 492 200 496 202
rect 492 199 493 200
rect 471 175 475 198
rect 478 198 493 199
rect 495 198 496 200
rect 478 195 496 198
rect 507 200 509 202
rect 511 200 512 202
rect 507 198 512 200
rect 541 205 542 207
rect 544 205 545 207
rect 478 190 482 195
rect 478 188 479 190
rect 481 188 482 190
rect 478 183 482 188
rect 478 179 486 183
rect 482 175 486 179
rect 471 174 478 175
rect 471 172 474 174
rect 476 172 478 174
rect 471 171 478 172
rect 482 174 499 175
rect 482 172 495 174
rect 497 172 499 174
rect 482 171 499 172
rect 507 174 511 198
rect 531 202 537 204
rect 541 203 545 205
rect 549 205 556 206
rect 549 203 552 205
rect 554 203 556 205
rect 531 200 532 202
rect 534 200 537 202
rect 531 198 537 200
rect 533 191 537 198
rect 549 202 556 203
rect 580 205 586 213
rect 618 211 620 213
rect 622 211 624 213
rect 618 210 624 211
rect 641 207 645 213
rect 580 203 582 205
rect 584 203 586 205
rect 580 202 586 203
rect 607 202 612 204
rect 533 190 546 191
rect 533 188 542 190
rect 544 188 546 190
rect 533 187 546 188
rect 533 183 537 187
rect 531 181 537 183
rect 531 179 532 181
rect 534 179 537 181
rect 531 177 537 179
rect 549 181 553 202
rect 549 179 550 181
rect 552 179 553 181
rect 549 177 553 179
rect 556 190 560 192
rect 556 188 557 190
rect 559 188 560 190
rect 556 174 560 188
rect 507 173 560 174
rect 507 171 509 173
rect 511 171 560 173
rect 507 170 560 171
rect 571 200 575 202
rect 571 198 572 200
rect 574 198 575 200
rect 592 200 596 202
rect 592 199 593 200
rect 571 175 575 198
rect 578 198 593 199
rect 595 198 596 200
rect 578 195 596 198
rect 607 200 609 202
rect 611 200 612 202
rect 607 198 612 200
rect 641 205 642 207
rect 644 205 645 207
rect 578 190 582 195
rect 578 188 579 190
rect 581 188 582 190
rect 578 183 582 188
rect 578 179 586 183
rect 582 175 586 179
rect 571 174 578 175
rect 571 172 574 174
rect 576 172 578 174
rect 571 171 578 172
rect 582 174 599 175
rect 582 172 595 174
rect 597 172 599 174
rect 582 171 599 172
rect 607 174 611 198
rect 631 202 637 204
rect 641 203 645 205
rect 649 205 656 206
rect 649 203 652 205
rect 654 203 656 205
rect 631 200 632 202
rect 634 200 637 202
rect 631 198 637 200
rect 633 191 637 198
rect 649 202 656 203
rect 680 205 686 213
rect 718 211 720 213
rect 722 211 724 213
rect 718 210 724 211
rect 741 207 745 213
rect 680 203 682 205
rect 684 203 686 205
rect 680 202 686 203
rect 707 202 712 204
rect 633 190 646 191
rect 633 188 642 190
rect 644 188 646 190
rect 633 187 646 188
rect 633 183 637 187
rect 631 181 637 183
rect 631 179 632 181
rect 634 179 637 181
rect 631 177 637 179
rect 649 181 653 202
rect 649 179 650 181
rect 652 179 653 181
rect 649 177 653 179
rect 656 190 660 192
rect 656 188 657 190
rect 659 188 660 190
rect 656 174 660 188
rect 607 173 660 174
rect 607 171 609 173
rect 611 171 660 173
rect 607 170 660 171
rect 671 200 675 202
rect 671 198 672 200
rect 674 198 675 200
rect 692 200 696 202
rect 692 199 693 200
rect 671 175 675 198
rect 678 198 693 199
rect 695 198 696 200
rect 678 195 696 198
rect 707 200 709 202
rect 711 200 712 202
rect 707 198 712 200
rect 741 205 742 207
rect 744 205 745 207
rect 678 190 682 195
rect 678 188 679 190
rect 681 188 682 190
rect 678 183 682 188
rect 678 179 686 183
rect 682 175 686 179
rect 671 174 678 175
rect 671 172 674 174
rect 676 172 678 174
rect 671 171 678 172
rect 682 174 699 175
rect 682 172 695 174
rect 697 172 699 174
rect 682 171 699 172
rect 707 174 711 198
rect 731 202 737 204
rect 741 203 745 205
rect 749 205 756 206
rect 749 203 752 205
rect 754 203 756 205
rect 731 200 732 202
rect 734 200 737 202
rect 731 198 737 200
rect 733 191 737 198
rect 749 202 756 203
rect 780 205 786 213
rect 780 203 782 205
rect 784 203 786 205
rect 780 202 786 203
rect 733 190 746 191
rect 733 188 742 190
rect 744 188 746 190
rect 733 187 746 188
rect 733 183 737 187
rect 731 181 737 183
rect 731 179 732 181
rect 734 179 737 181
rect 731 177 737 179
rect 749 181 753 202
rect 749 179 750 181
rect 752 179 753 181
rect 749 177 753 179
rect 756 190 760 192
rect 756 188 757 190
rect 759 188 760 190
rect 756 174 760 188
rect 707 173 760 174
rect 707 171 709 173
rect 711 171 760 173
rect 707 170 760 171
rect 771 200 775 202
rect 771 198 772 200
rect 774 198 775 200
rect 792 200 796 202
rect 792 199 793 200
rect 771 175 775 198
rect 778 198 793 199
rect 795 198 796 200
rect 778 195 796 198
rect 778 190 782 195
rect 778 188 779 190
rect 781 188 782 190
rect 778 183 782 188
rect 778 179 786 183
rect 782 175 786 179
rect 771 174 778 175
rect 771 172 774 174
rect 776 172 778 174
rect 771 171 778 172
rect 782 174 799 175
rect 782 172 795 174
rect 797 172 799 174
rect 782 171 799 172
rect 17 165 23 166
rect 17 163 19 165
rect 21 163 23 165
rect 17 157 23 163
rect 36 165 42 166
rect 36 163 38 165
rect 40 163 42 165
rect 80 166 86 167
rect 80 164 82 166
rect 84 164 86 166
rect 36 157 42 163
rect 80 157 86 164
rect 117 165 123 166
rect 117 163 119 165
rect 121 163 123 165
rect 117 157 123 163
rect 136 165 142 166
rect 136 163 138 165
rect 140 163 142 165
rect 180 166 186 167
rect 180 164 182 166
rect 184 164 186 166
rect 136 157 142 163
rect 180 157 186 164
rect 217 165 223 166
rect 217 163 219 165
rect 221 163 223 165
rect 217 157 223 163
rect 236 165 242 166
rect 236 163 238 165
rect 240 163 242 165
rect 280 166 286 167
rect 280 164 282 166
rect 284 164 286 166
rect 236 157 242 163
rect 280 157 286 164
rect 317 165 323 166
rect 317 163 319 165
rect 321 163 323 165
rect 317 157 323 163
rect 336 165 342 166
rect 336 163 338 165
rect 340 163 342 165
rect 380 166 386 167
rect 380 164 382 166
rect 384 164 386 166
rect 336 157 342 163
rect 380 157 386 164
rect 419 165 425 166
rect 419 163 421 165
rect 423 163 425 165
rect 419 157 425 163
rect 438 165 444 166
rect 438 163 440 165
rect 442 163 444 165
rect 482 166 488 167
rect 482 164 484 166
rect 486 164 488 166
rect 438 157 444 163
rect 482 157 488 164
rect 519 165 525 166
rect 519 163 521 165
rect 523 163 525 165
rect 519 157 525 163
rect 538 165 544 166
rect 538 163 540 165
rect 542 163 544 165
rect 582 166 588 167
rect 582 164 584 166
rect 586 164 588 166
rect 538 157 544 163
rect 582 157 588 164
rect 619 165 625 166
rect 619 163 621 165
rect 623 163 625 165
rect 619 157 625 163
rect 638 165 644 166
rect 638 163 640 165
rect 642 163 644 165
rect 682 166 688 167
rect 682 164 684 166
rect 686 164 688 166
rect 638 157 644 163
rect 682 157 688 164
rect 719 165 725 166
rect 719 163 721 165
rect 723 163 725 165
rect 719 157 725 163
rect 738 165 744 166
rect 738 163 740 165
rect 742 163 744 165
rect 782 166 788 167
rect 782 164 784 166
rect 786 164 788 166
rect 738 157 744 163
rect 782 157 788 164
rect 17 135 23 141
rect 17 133 19 135
rect 21 133 23 135
rect 17 132 23 133
rect 36 135 42 141
rect 36 133 38 135
rect 40 133 42 135
rect 36 132 42 133
rect 80 134 86 141
rect 80 132 82 134
rect 84 132 86 134
rect 117 135 123 141
rect 117 133 119 135
rect 121 133 123 135
rect 117 132 123 133
rect 136 135 142 141
rect 136 133 138 135
rect 140 133 142 135
rect 136 132 142 133
rect 80 131 86 132
rect 180 134 186 141
rect 180 132 182 134
rect 184 132 186 134
rect 217 135 223 141
rect 217 133 219 135
rect 221 133 223 135
rect 217 132 223 133
rect 236 135 242 141
rect 236 133 238 135
rect 240 133 242 135
rect 236 132 242 133
rect 180 131 186 132
rect 280 134 286 141
rect 280 132 282 134
rect 284 132 286 134
rect 317 135 323 141
rect 317 133 319 135
rect 321 133 323 135
rect 317 132 323 133
rect 336 135 342 141
rect 336 133 338 135
rect 340 133 342 135
rect 336 132 342 133
rect 280 131 286 132
rect 380 134 386 141
rect 380 132 382 134
rect 384 132 386 134
rect 419 135 425 141
rect 419 133 421 135
rect 423 133 425 135
rect 419 132 425 133
rect 438 135 444 141
rect 438 133 440 135
rect 442 133 444 135
rect 438 132 444 133
rect 380 131 386 132
rect 482 134 488 141
rect 482 132 484 134
rect 486 132 488 134
rect 519 135 525 141
rect 519 133 521 135
rect 523 133 525 135
rect 519 132 525 133
rect 538 135 544 141
rect 538 133 540 135
rect 542 133 544 135
rect 538 132 544 133
rect 482 131 488 132
rect 582 134 588 141
rect 582 132 584 134
rect 586 132 588 134
rect 619 135 625 141
rect 619 133 621 135
rect 623 133 625 135
rect 619 132 625 133
rect 638 135 644 141
rect 638 133 640 135
rect 642 133 644 135
rect 638 132 644 133
rect 582 131 588 132
rect 682 134 688 141
rect 682 132 684 134
rect 686 132 688 134
rect 719 135 725 141
rect 719 133 721 135
rect 723 133 725 135
rect 719 132 725 133
rect 738 135 744 141
rect 738 133 740 135
rect 742 133 744 135
rect 738 132 744 133
rect 682 131 688 132
rect 782 134 788 141
rect 782 132 784 134
rect 786 132 788 134
rect 782 131 788 132
rect 5 127 58 128
rect 5 125 7 127
rect 9 125 58 127
rect 5 124 58 125
rect 5 100 9 124
rect 29 119 35 121
rect 29 117 30 119
rect 32 117 35 119
rect 29 115 35 117
rect 31 111 35 115
rect 47 119 51 121
rect 47 117 48 119
rect 50 117 51 119
rect 31 110 44 111
rect 31 108 40 110
rect 42 108 44 110
rect 31 107 44 108
rect 5 98 10 100
rect 5 96 7 98
rect 9 96 10 98
rect 5 94 10 96
rect 31 100 35 107
rect 29 98 35 100
rect 29 96 30 98
rect 32 96 35 98
rect 29 94 35 96
rect 47 96 51 117
rect 54 110 58 124
rect 54 108 55 110
rect 57 108 58 110
rect 54 106 58 108
rect 105 127 158 128
rect 69 126 76 127
rect 69 124 72 126
rect 74 124 76 126
rect 69 123 76 124
rect 80 126 97 127
rect 80 124 93 126
rect 95 124 97 126
rect 80 123 97 124
rect 105 125 107 127
rect 109 125 158 127
rect 105 124 158 125
rect 69 100 73 123
rect 80 119 84 123
rect 69 98 70 100
rect 72 98 73 100
rect 76 115 84 119
rect 76 110 80 115
rect 76 108 77 110
rect 79 108 80 110
rect 76 103 80 108
rect 76 100 94 103
rect 76 99 91 100
rect 69 96 73 98
rect 90 98 91 99
rect 93 98 94 100
rect 90 96 94 98
rect 105 100 109 124
rect 129 119 135 121
rect 129 117 130 119
rect 132 117 135 119
rect 129 115 135 117
rect 131 111 135 115
rect 147 119 151 121
rect 147 117 148 119
rect 150 117 151 119
rect 131 110 144 111
rect 131 108 140 110
rect 142 108 144 110
rect 131 107 144 108
rect 105 98 110 100
rect 105 96 107 98
rect 109 96 110 98
rect 47 95 54 96
rect 39 93 43 95
rect 39 91 40 93
rect 42 91 43 93
rect 47 93 50 95
rect 52 93 54 95
rect 47 92 54 93
rect 78 95 84 96
rect 78 93 80 95
rect 82 93 84 95
rect 105 94 110 96
rect 131 100 135 107
rect 129 98 135 100
rect 129 96 130 98
rect 132 96 135 98
rect 129 94 135 96
rect 147 96 151 117
rect 154 110 158 124
rect 154 108 155 110
rect 157 108 158 110
rect 154 106 158 108
rect 205 127 258 128
rect 169 126 176 127
rect 169 124 172 126
rect 174 124 176 126
rect 169 123 176 124
rect 180 126 197 127
rect 180 124 193 126
rect 195 124 197 126
rect 180 123 197 124
rect 205 125 207 127
rect 209 125 258 127
rect 205 124 258 125
rect 169 100 173 123
rect 180 119 184 123
rect 169 98 170 100
rect 172 98 173 100
rect 176 115 184 119
rect 176 110 180 115
rect 176 108 177 110
rect 179 108 180 110
rect 176 103 180 108
rect 176 100 194 103
rect 176 99 191 100
rect 169 96 173 98
rect 190 98 191 99
rect 193 98 194 100
rect 190 96 194 98
rect 205 100 209 124
rect 229 119 235 121
rect 229 117 230 119
rect 232 117 235 119
rect 229 115 235 117
rect 231 111 235 115
rect 247 119 251 121
rect 247 117 248 119
rect 250 117 251 119
rect 231 110 244 111
rect 205 98 210 100
rect 205 96 207 98
rect 209 96 210 98
rect 147 95 154 96
rect 16 87 22 88
rect 16 85 18 87
rect 20 85 22 87
rect 39 85 43 91
rect 78 85 84 93
rect 139 93 143 95
rect 139 91 140 93
rect 142 91 143 93
rect 147 93 150 95
rect 152 93 154 95
rect 147 92 154 93
rect 178 95 184 96
rect 178 93 180 95
rect 182 93 184 95
rect 205 94 210 96
rect 231 108 240 110
rect 242 108 244 110
rect 231 107 244 108
rect 231 100 235 107
rect 229 98 235 100
rect 229 96 230 98
rect 232 96 235 98
rect 229 94 235 96
rect 247 96 251 117
rect 254 110 258 124
rect 254 108 255 110
rect 257 108 258 110
rect 254 106 258 108
rect 305 127 358 128
rect 269 126 276 127
rect 269 124 272 126
rect 274 124 276 126
rect 269 123 276 124
rect 280 126 297 127
rect 280 124 293 126
rect 295 124 297 126
rect 280 123 297 124
rect 305 125 307 127
rect 309 125 358 127
rect 305 124 358 125
rect 269 100 273 123
rect 280 119 284 123
rect 269 98 270 100
rect 272 98 273 100
rect 276 115 284 119
rect 276 110 280 115
rect 276 108 277 110
rect 279 108 280 110
rect 276 103 280 108
rect 276 100 294 103
rect 276 99 291 100
rect 269 96 273 98
rect 290 98 291 99
rect 293 98 294 100
rect 290 96 294 98
rect 305 100 309 124
rect 329 119 335 121
rect 329 117 330 119
rect 332 117 335 119
rect 329 115 335 117
rect 331 111 335 115
rect 347 119 351 121
rect 347 117 348 119
rect 350 117 351 119
rect 331 110 344 111
rect 331 108 340 110
rect 342 108 344 110
rect 331 107 344 108
rect 305 98 310 100
rect 305 96 307 98
rect 309 96 310 98
rect 247 95 254 96
rect 116 87 122 88
rect 116 85 118 87
rect 120 85 122 87
rect 139 85 143 91
rect 178 85 184 93
rect 239 93 243 95
rect 239 91 240 93
rect 242 91 243 93
rect 247 93 250 95
rect 252 93 254 95
rect 247 92 254 93
rect 278 95 284 96
rect 278 93 280 95
rect 282 93 284 95
rect 305 94 310 96
rect 331 100 335 107
rect 329 98 335 100
rect 329 96 330 98
rect 332 96 335 98
rect 329 94 335 96
rect 347 96 351 117
rect 354 110 358 124
rect 354 108 355 110
rect 357 108 358 110
rect 354 106 358 108
rect 407 127 460 128
rect 369 126 376 127
rect 369 124 372 126
rect 374 124 376 126
rect 369 123 376 124
rect 380 126 397 127
rect 380 124 393 126
rect 395 124 397 126
rect 380 123 397 124
rect 407 125 409 127
rect 411 125 460 127
rect 407 124 460 125
rect 369 100 373 123
rect 380 119 384 123
rect 369 98 370 100
rect 372 98 373 100
rect 376 115 384 119
rect 376 110 380 115
rect 376 108 377 110
rect 379 108 380 110
rect 376 103 380 108
rect 376 100 394 103
rect 376 99 391 100
rect 369 96 373 98
rect 390 98 391 99
rect 393 98 394 100
rect 390 96 394 98
rect 407 100 411 124
rect 431 119 437 121
rect 431 117 432 119
rect 434 117 437 119
rect 431 115 437 117
rect 433 111 437 115
rect 449 119 453 121
rect 449 117 450 119
rect 452 117 453 119
rect 433 110 446 111
rect 433 108 442 110
rect 444 108 446 110
rect 433 107 446 108
rect 407 98 412 100
rect 407 96 409 98
rect 411 96 412 98
rect 347 95 354 96
rect 216 87 222 88
rect 216 85 218 87
rect 220 85 222 87
rect 239 85 243 91
rect 278 85 284 93
rect 339 93 343 95
rect 339 91 340 93
rect 342 91 343 93
rect 347 93 350 95
rect 352 93 354 95
rect 347 92 354 93
rect 378 95 384 96
rect 378 93 380 95
rect 382 93 384 95
rect 407 94 412 96
rect 433 100 437 107
rect 431 98 437 100
rect 431 96 432 98
rect 434 96 437 98
rect 431 94 437 96
rect 449 96 453 117
rect 456 110 460 124
rect 456 108 457 110
rect 459 108 460 110
rect 456 106 460 108
rect 507 127 560 128
rect 471 126 478 127
rect 471 124 474 126
rect 476 124 478 126
rect 471 123 478 124
rect 482 126 499 127
rect 482 124 495 126
rect 497 124 499 126
rect 482 123 499 124
rect 507 125 509 127
rect 511 125 560 127
rect 507 124 560 125
rect 471 100 475 123
rect 482 119 486 123
rect 471 98 472 100
rect 474 98 475 100
rect 478 115 486 119
rect 478 110 482 115
rect 478 108 479 110
rect 481 108 482 110
rect 478 103 482 108
rect 478 100 496 103
rect 478 99 493 100
rect 471 96 475 98
rect 492 98 493 99
rect 495 98 496 100
rect 492 96 496 98
rect 507 100 511 124
rect 531 119 537 121
rect 531 117 532 119
rect 534 117 537 119
rect 531 115 537 117
rect 533 111 537 115
rect 549 119 553 121
rect 549 117 550 119
rect 552 117 553 119
rect 533 110 546 111
rect 533 108 542 110
rect 544 108 546 110
rect 533 107 546 108
rect 507 98 512 100
rect 507 96 509 98
rect 511 96 512 98
rect 449 95 456 96
rect 316 87 322 88
rect 316 85 318 87
rect 320 85 322 87
rect 339 85 343 91
rect 378 85 384 93
rect 441 93 445 95
rect 441 91 442 93
rect 444 91 445 93
rect 449 93 452 95
rect 454 93 456 95
rect 449 92 456 93
rect 480 95 486 96
rect 480 93 482 95
rect 484 93 486 95
rect 507 94 512 96
rect 533 100 537 107
rect 531 98 537 100
rect 531 96 532 98
rect 534 96 537 98
rect 531 94 537 96
rect 549 96 553 117
rect 556 110 560 124
rect 556 108 557 110
rect 559 108 560 110
rect 556 106 560 108
rect 607 127 660 128
rect 571 126 578 127
rect 571 124 574 126
rect 576 124 578 126
rect 571 123 578 124
rect 582 126 599 127
rect 582 124 595 126
rect 597 124 599 126
rect 582 123 599 124
rect 607 125 609 127
rect 611 125 660 127
rect 607 124 660 125
rect 571 100 575 123
rect 582 119 586 123
rect 571 98 572 100
rect 574 98 575 100
rect 578 115 586 119
rect 578 110 582 115
rect 578 108 579 110
rect 581 108 582 110
rect 578 103 582 108
rect 578 100 596 103
rect 607 100 611 124
rect 631 119 637 121
rect 631 117 632 119
rect 634 117 637 119
rect 631 115 637 117
rect 633 111 637 115
rect 649 119 653 121
rect 649 117 650 119
rect 652 117 653 119
rect 633 110 646 111
rect 633 108 642 110
rect 644 108 646 110
rect 633 107 646 108
rect 578 99 593 100
rect 571 96 575 98
rect 592 98 593 99
rect 595 98 596 100
rect 592 96 596 98
rect 607 98 612 100
rect 607 96 609 98
rect 611 96 612 98
rect 549 95 556 96
rect 418 87 424 88
rect 418 85 420 87
rect 422 85 424 87
rect 441 85 445 91
rect 480 85 486 93
rect 541 93 545 95
rect 541 91 542 93
rect 544 91 545 93
rect 549 93 552 95
rect 554 93 556 95
rect 549 92 556 93
rect 580 95 586 96
rect 580 93 582 95
rect 584 93 586 95
rect 607 94 612 96
rect 633 100 637 107
rect 631 98 637 100
rect 631 96 632 98
rect 634 96 637 98
rect 631 94 637 96
rect 649 96 653 117
rect 656 110 660 124
rect 656 108 657 110
rect 659 108 660 110
rect 656 106 660 108
rect 707 127 760 128
rect 671 126 678 127
rect 671 124 674 126
rect 676 124 678 126
rect 671 123 678 124
rect 682 126 699 127
rect 682 124 695 126
rect 697 124 699 126
rect 682 123 699 124
rect 707 125 709 127
rect 711 125 760 127
rect 707 124 760 125
rect 671 100 675 123
rect 682 119 686 123
rect 671 98 672 100
rect 674 98 675 100
rect 678 115 686 119
rect 678 110 682 115
rect 678 108 679 110
rect 681 108 682 110
rect 678 103 682 108
rect 678 100 696 103
rect 678 99 693 100
rect 671 96 675 98
rect 692 98 693 99
rect 695 98 696 100
rect 692 96 696 98
rect 707 100 711 124
rect 731 119 737 121
rect 731 117 732 119
rect 734 117 737 119
rect 731 115 737 117
rect 733 111 737 115
rect 749 119 753 121
rect 749 117 750 119
rect 752 117 753 119
rect 733 110 746 111
rect 707 98 712 100
rect 707 96 709 98
rect 711 96 712 98
rect 649 95 656 96
rect 518 87 524 88
rect 518 85 520 87
rect 522 85 524 87
rect 541 85 545 91
rect 580 85 586 93
rect 641 93 645 95
rect 641 91 642 93
rect 644 91 645 93
rect 649 93 652 95
rect 654 93 656 95
rect 649 92 656 93
rect 680 95 686 96
rect 680 93 682 95
rect 684 93 686 95
rect 707 94 712 96
rect 733 108 742 110
rect 744 108 746 110
rect 733 107 746 108
rect 733 100 737 107
rect 731 98 737 100
rect 731 96 732 98
rect 734 96 737 98
rect 731 94 737 96
rect 749 96 753 117
rect 756 110 760 124
rect 756 108 757 110
rect 759 108 760 110
rect 756 106 760 108
rect 771 126 778 127
rect 771 124 774 126
rect 776 124 778 126
rect 771 123 778 124
rect 782 126 799 127
rect 782 124 795 126
rect 797 124 799 126
rect 782 123 799 124
rect 771 100 775 123
rect 782 119 786 123
rect 771 98 772 100
rect 774 98 775 100
rect 778 115 786 119
rect 778 110 782 115
rect 778 108 779 110
rect 781 108 782 110
rect 778 103 782 108
rect 778 100 796 103
rect 778 99 793 100
rect 771 96 775 98
rect 792 98 793 99
rect 795 98 796 100
rect 792 96 796 98
rect 749 95 756 96
rect 618 87 624 88
rect 618 85 620 87
rect 622 85 624 87
rect 641 85 645 91
rect 680 85 686 93
rect 741 93 745 95
rect 741 91 742 93
rect 744 91 745 93
rect 749 93 752 95
rect 754 93 756 95
rect 749 92 756 93
rect 780 95 786 96
rect 780 93 782 95
rect 784 93 786 95
rect 718 87 724 88
rect 718 85 720 87
rect 722 85 724 87
rect 741 85 745 91
rect 780 85 786 93
rect 18 61 24 69
rect 59 63 63 69
rect 81 67 82 69
rect 84 67 86 69
rect 81 66 86 67
rect 18 59 20 61
rect 22 59 24 61
rect 18 58 24 59
rect 48 61 55 62
rect 48 59 50 61
rect 52 59 55 61
rect 59 61 60 63
rect 62 61 63 63
rect 59 59 63 61
rect 48 58 55 59
rect 8 56 12 58
rect 8 54 9 56
rect 11 55 12 56
rect 29 56 33 58
rect 11 54 26 55
rect 8 51 26 54
rect 22 46 26 51
rect 22 44 23 46
rect 25 44 26 46
rect 22 39 26 44
rect 18 35 26 39
rect 29 54 30 56
rect 32 54 33 56
rect 18 31 22 35
rect 29 31 33 54
rect 5 30 22 31
rect 5 28 7 30
rect 9 28 22 30
rect 5 27 22 28
rect 26 30 33 31
rect 26 28 28 30
rect 30 28 33 30
rect 26 27 33 28
rect 44 46 48 48
rect 44 44 45 46
rect 47 44 48 46
rect 44 30 48 44
rect 51 37 55 58
rect 67 58 73 60
rect 67 56 70 58
rect 72 56 73 58
rect 67 54 73 56
rect 67 47 71 54
rect 58 46 71 47
rect 58 44 60 46
rect 62 44 71 46
rect 118 61 124 69
rect 159 63 163 69
rect 180 67 182 69
rect 184 67 186 69
rect 180 66 186 67
rect 92 58 97 60
rect 118 59 120 61
rect 122 59 124 61
rect 118 58 124 59
rect 148 61 155 62
rect 148 59 150 61
rect 152 59 155 61
rect 159 61 160 63
rect 162 61 163 63
rect 159 59 163 61
rect 148 58 155 59
rect 92 56 93 58
rect 95 56 97 58
rect 92 54 97 56
rect 58 43 71 44
rect 51 35 52 37
rect 54 35 55 37
rect 51 33 55 35
rect 67 39 71 43
rect 67 37 73 39
rect 67 35 70 37
rect 72 35 73 37
rect 67 33 73 35
rect 93 30 97 54
rect 108 56 112 58
rect 108 54 109 56
rect 111 55 112 56
rect 129 56 133 58
rect 111 54 126 55
rect 108 51 126 54
rect 122 46 126 51
rect 122 44 123 46
rect 125 44 126 46
rect 122 39 126 44
rect 118 35 126 39
rect 129 54 130 56
rect 132 54 133 56
rect 118 31 122 35
rect 129 31 133 54
rect 44 29 97 30
rect 44 27 93 29
rect 95 27 97 29
rect 109 27 122 31
rect 126 30 133 31
rect 126 28 128 30
rect 130 28 133 30
rect 126 27 133 28
rect 44 26 97 27
rect 144 46 148 48
rect 144 44 145 46
rect 147 44 148 46
rect 144 30 148 44
rect 151 37 155 58
rect 167 58 173 60
rect 167 56 170 58
rect 172 56 173 58
rect 167 54 173 56
rect 167 47 171 54
rect 158 46 171 47
rect 158 44 160 46
rect 162 44 171 46
rect 218 61 224 69
rect 259 63 263 69
rect 280 67 282 69
rect 284 67 286 69
rect 280 66 286 67
rect 192 58 197 60
rect 218 59 220 61
rect 222 59 224 61
rect 218 58 224 59
rect 248 61 255 62
rect 248 59 250 61
rect 252 59 255 61
rect 259 61 260 63
rect 262 61 263 63
rect 259 59 263 61
rect 248 58 255 59
rect 192 56 193 58
rect 195 56 197 58
rect 192 54 197 56
rect 158 43 171 44
rect 151 35 152 37
rect 154 35 155 37
rect 151 33 155 35
rect 167 39 171 43
rect 167 37 173 39
rect 167 35 170 37
rect 172 35 173 37
rect 167 33 173 35
rect 193 30 197 54
rect 208 56 212 58
rect 208 54 209 56
rect 211 55 212 56
rect 229 56 233 58
rect 211 54 226 55
rect 208 51 226 54
rect 222 46 226 51
rect 222 44 223 46
rect 225 44 226 46
rect 222 39 226 44
rect 218 35 226 39
rect 229 54 230 56
rect 232 54 233 56
rect 218 31 222 35
rect 229 31 233 54
rect 144 29 197 30
rect 144 27 193 29
rect 195 27 197 29
rect 205 30 222 31
rect 205 28 207 30
rect 209 28 222 30
rect 205 27 222 28
rect 226 30 233 31
rect 226 28 228 30
rect 230 28 233 30
rect 226 27 233 28
rect 144 26 197 27
rect 244 46 248 48
rect 244 44 245 46
rect 247 44 248 46
rect 244 30 248 44
rect 251 37 255 58
rect 267 58 273 60
rect 267 56 270 58
rect 272 56 273 58
rect 267 54 273 56
rect 267 47 271 54
rect 258 46 271 47
rect 258 44 260 46
rect 262 44 271 46
rect 318 61 324 69
rect 359 63 363 69
rect 380 67 382 69
rect 384 67 386 69
rect 380 66 386 67
rect 292 58 297 60
rect 318 59 320 61
rect 322 59 324 61
rect 318 58 324 59
rect 348 61 355 62
rect 348 59 350 61
rect 352 59 355 61
rect 359 61 360 63
rect 362 61 363 63
rect 359 59 363 61
rect 348 58 355 59
rect 292 56 293 58
rect 295 56 297 58
rect 292 54 297 56
rect 258 43 271 44
rect 251 35 252 37
rect 254 35 255 37
rect 251 33 255 35
rect 267 39 271 43
rect 267 37 273 39
rect 267 35 270 37
rect 272 35 273 37
rect 267 33 273 35
rect 293 30 297 54
rect 308 56 312 58
rect 308 54 309 56
rect 311 55 312 56
rect 329 56 333 58
rect 311 54 326 55
rect 308 51 326 54
rect 322 46 326 51
rect 322 44 323 46
rect 325 44 326 46
rect 322 39 326 44
rect 318 35 326 39
rect 329 54 330 56
rect 332 54 333 56
rect 318 31 322 35
rect 329 31 333 54
rect 244 29 297 30
rect 244 27 293 29
rect 295 27 297 29
rect 305 30 322 31
rect 305 28 307 30
rect 309 28 322 30
rect 305 27 322 28
rect 326 30 333 31
rect 326 28 328 30
rect 330 28 333 30
rect 326 27 333 28
rect 244 26 297 27
rect 344 46 348 48
rect 344 44 345 46
rect 347 44 348 46
rect 344 30 348 44
rect 351 37 355 58
rect 367 58 373 60
rect 418 61 424 69
rect 459 63 463 69
rect 480 67 482 69
rect 484 67 486 69
rect 480 66 486 67
rect 367 56 370 58
rect 372 56 373 58
rect 367 54 373 56
rect 367 47 371 54
rect 392 58 397 60
rect 418 59 420 61
rect 422 59 424 61
rect 418 58 424 59
rect 448 61 455 62
rect 448 59 450 61
rect 452 59 455 61
rect 459 61 460 63
rect 462 61 463 63
rect 459 59 463 61
rect 448 58 455 59
rect 392 56 393 58
rect 395 56 397 58
rect 392 54 397 56
rect 358 46 371 47
rect 358 44 360 46
rect 362 44 371 46
rect 358 43 371 44
rect 351 35 352 37
rect 354 35 355 37
rect 351 33 355 35
rect 367 39 371 43
rect 367 37 373 39
rect 367 35 370 37
rect 372 35 373 37
rect 367 33 373 35
rect 393 30 397 54
rect 408 56 412 58
rect 408 54 409 56
rect 411 55 412 56
rect 429 56 433 58
rect 411 54 426 55
rect 408 51 426 54
rect 422 46 426 51
rect 422 44 423 46
rect 425 44 426 46
rect 422 39 426 44
rect 418 35 426 39
rect 429 54 430 56
rect 432 54 433 56
rect 418 31 422 35
rect 429 31 433 54
rect 344 29 397 30
rect 344 27 393 29
rect 395 27 397 29
rect 405 30 422 31
rect 405 28 407 30
rect 409 28 422 30
rect 405 27 422 28
rect 426 30 433 31
rect 426 28 428 30
rect 430 28 433 30
rect 426 27 433 28
rect 344 26 397 27
rect 444 46 448 48
rect 444 44 445 46
rect 447 44 448 46
rect 444 30 448 44
rect 451 37 455 58
rect 467 58 473 60
rect 467 56 470 58
rect 472 56 473 58
rect 467 54 473 56
rect 467 47 471 54
rect 492 58 497 60
rect 492 56 493 58
rect 495 56 497 58
rect 492 54 497 56
rect 458 46 471 47
rect 458 44 460 46
rect 462 44 471 46
rect 458 43 471 44
rect 451 35 452 37
rect 454 35 455 37
rect 451 33 455 35
rect 467 39 471 43
rect 467 37 473 39
rect 467 35 470 37
rect 472 35 473 37
rect 467 33 473 35
rect 493 30 497 54
rect 518 61 524 69
rect 559 63 563 69
rect 580 67 582 69
rect 584 67 586 69
rect 580 66 586 67
rect 518 59 520 61
rect 522 59 524 61
rect 518 58 524 59
rect 548 61 555 62
rect 548 59 550 61
rect 552 59 555 61
rect 559 61 560 63
rect 562 61 563 63
rect 559 59 563 61
rect 548 58 555 59
rect 508 56 512 58
rect 508 54 509 56
rect 511 55 512 56
rect 529 56 533 58
rect 511 54 526 55
rect 508 51 526 54
rect 522 46 526 51
rect 522 44 523 46
rect 525 44 526 46
rect 522 39 526 44
rect 518 35 526 39
rect 529 54 530 56
rect 532 54 533 56
rect 518 31 522 35
rect 529 31 533 54
rect 444 29 497 30
rect 444 27 493 29
rect 495 27 497 29
rect 505 30 522 31
rect 505 28 507 30
rect 509 28 522 30
rect 505 27 522 28
rect 526 30 533 31
rect 526 28 528 30
rect 530 28 533 30
rect 526 27 533 28
rect 444 26 497 27
rect 544 46 548 48
rect 544 44 545 46
rect 547 44 548 46
rect 544 30 548 44
rect 551 37 555 58
rect 567 58 573 60
rect 567 56 570 58
rect 572 56 573 58
rect 567 54 573 56
rect 567 47 571 54
rect 592 58 597 60
rect 592 56 593 58
rect 595 56 597 58
rect 592 54 597 56
rect 558 46 571 47
rect 558 44 560 46
rect 562 44 571 46
rect 558 43 571 44
rect 551 35 552 37
rect 554 35 555 37
rect 551 33 555 35
rect 567 39 571 43
rect 567 37 573 39
rect 567 35 570 37
rect 572 35 573 37
rect 567 33 573 35
rect 593 30 597 54
rect 618 61 624 69
rect 659 63 663 69
rect 680 67 682 69
rect 684 67 686 69
rect 680 66 686 67
rect 618 59 620 61
rect 622 59 624 61
rect 618 58 624 59
rect 648 61 655 62
rect 648 59 650 61
rect 652 59 655 61
rect 659 61 660 63
rect 662 61 663 63
rect 659 59 663 61
rect 648 58 655 59
rect 608 56 612 58
rect 608 54 609 56
rect 611 55 612 56
rect 629 56 633 58
rect 611 54 626 55
rect 608 51 626 54
rect 622 46 626 51
rect 622 44 623 46
rect 625 44 626 46
rect 622 39 626 44
rect 618 35 626 39
rect 629 54 630 56
rect 632 54 633 56
rect 618 31 622 35
rect 629 31 633 54
rect 544 29 597 30
rect 544 27 593 29
rect 595 27 597 29
rect 605 30 622 31
rect 605 28 607 30
rect 609 28 622 30
rect 605 27 622 28
rect 626 30 633 31
rect 626 28 628 30
rect 630 28 633 30
rect 626 27 633 28
rect 544 26 597 27
rect 644 46 648 48
rect 644 44 645 46
rect 647 44 648 46
rect 644 30 648 44
rect 651 37 655 58
rect 667 58 673 60
rect 667 56 670 58
rect 672 56 673 58
rect 667 54 673 56
rect 667 47 671 54
rect 692 58 697 60
rect 692 56 693 58
rect 695 56 697 58
rect 692 54 697 56
rect 658 46 671 47
rect 658 44 660 46
rect 662 44 671 46
rect 658 43 671 44
rect 651 35 652 37
rect 654 35 655 37
rect 651 33 655 35
rect 667 39 671 43
rect 667 37 673 39
rect 667 35 670 37
rect 672 35 673 37
rect 667 33 673 35
rect 693 30 697 54
rect 718 61 724 69
rect 759 63 763 69
rect 780 67 782 69
rect 784 67 786 69
rect 780 66 786 67
rect 718 59 720 61
rect 722 59 724 61
rect 718 58 724 59
rect 748 61 755 62
rect 748 59 750 61
rect 752 59 755 61
rect 759 61 760 63
rect 762 61 763 63
rect 759 59 763 61
rect 748 58 755 59
rect 708 56 712 58
rect 708 54 709 56
rect 711 55 712 56
rect 729 56 733 58
rect 711 54 726 55
rect 708 51 726 54
rect 722 46 726 51
rect 722 44 723 46
rect 725 44 726 46
rect 722 39 726 44
rect 718 35 726 39
rect 729 54 730 56
rect 732 54 733 56
rect 718 31 722 35
rect 729 31 733 54
rect 644 29 697 30
rect 644 27 693 29
rect 695 27 697 29
rect 705 30 722 31
rect 705 28 707 30
rect 709 28 722 30
rect 705 27 722 28
rect 726 30 733 31
rect 726 28 728 30
rect 730 28 733 30
rect 726 27 733 28
rect 644 26 697 27
rect 744 46 748 48
rect 744 44 745 46
rect 747 44 748 46
rect 744 30 748 44
rect 751 37 755 58
rect 767 58 773 60
rect 767 56 770 58
rect 772 56 773 58
rect 767 54 773 56
rect 767 47 771 54
rect 792 58 797 60
rect 792 56 793 58
rect 795 56 797 58
rect 792 54 797 56
rect 758 46 771 47
rect 758 44 760 46
rect 762 44 771 46
rect 758 43 771 44
rect 751 35 752 37
rect 754 35 755 37
rect 751 33 755 35
rect 767 39 771 43
rect 767 37 773 39
rect 767 35 770 37
rect 772 35 773 37
rect 767 33 773 35
rect 793 30 797 54
rect 744 29 797 30
rect 744 27 793 29
rect 795 27 797 29
rect 744 26 797 27
rect 16 22 22 23
rect 16 20 18 22
rect 20 20 22 22
rect 16 13 22 20
rect 116 22 122 23
rect 60 21 66 22
rect 60 19 62 21
rect 64 19 66 21
rect 60 13 66 19
rect 79 21 85 22
rect 79 19 81 21
rect 83 19 85 21
rect 79 13 85 19
rect 116 20 118 22
rect 120 20 122 22
rect 116 13 122 20
rect 216 22 222 23
rect 160 21 166 22
rect 160 19 162 21
rect 164 19 166 21
rect 160 13 166 19
rect 179 21 185 22
rect 179 19 181 21
rect 183 19 185 21
rect 179 13 185 19
rect 216 20 218 22
rect 220 20 222 22
rect 216 13 222 20
rect 316 22 322 23
rect 260 21 266 22
rect 260 19 262 21
rect 264 19 266 21
rect 260 13 266 19
rect 279 21 285 22
rect 279 19 281 21
rect 283 19 285 21
rect 279 13 285 19
rect 316 20 318 22
rect 320 20 322 22
rect 316 13 322 20
rect 416 22 422 23
rect 360 21 366 22
rect 360 19 362 21
rect 364 19 366 21
rect 360 13 366 19
rect 379 21 385 22
rect 379 19 381 21
rect 383 19 385 21
rect 379 13 385 19
rect 416 20 418 22
rect 420 20 422 22
rect 416 13 422 20
rect 516 22 522 23
rect 460 21 466 22
rect 460 19 462 21
rect 464 19 466 21
rect 460 13 466 19
rect 479 21 485 22
rect 479 19 481 21
rect 483 19 485 21
rect 479 13 485 19
rect 516 20 518 22
rect 520 20 522 22
rect 516 13 522 20
rect 616 22 622 23
rect 560 21 566 22
rect 560 19 562 21
rect 564 19 566 21
rect 560 13 566 19
rect 579 21 585 22
rect 579 19 581 21
rect 583 19 585 21
rect 579 13 585 19
rect 616 20 618 22
rect 620 20 622 22
rect 616 13 622 20
rect 716 22 722 23
rect 660 21 666 22
rect 660 19 662 21
rect 664 19 666 21
rect 660 13 666 19
rect 679 21 685 22
rect 679 19 681 21
rect 683 19 685 21
rect 679 13 685 19
rect 716 20 718 22
rect 720 20 722 22
rect 716 13 722 20
rect 760 21 766 22
rect 760 19 762 21
rect 764 19 766 21
rect 760 13 766 19
rect 779 21 785 22
rect 779 19 781 21
rect 783 19 785 21
rect 779 13 785 19
rect -1 -38 5 -31
rect 43 -37 49 -31
rect -1 -40 1 -38
rect 3 -40 5 -38
rect -1 -41 5 -40
rect 43 -39 45 -37
rect 47 -39 49 -37
rect 43 -40 49 -39
rect 62 -37 68 -31
rect 62 -39 64 -37
rect 66 -39 68 -37
rect 62 -40 68 -39
rect 105 -38 111 -31
rect 149 -37 155 -31
rect 105 -40 107 -38
rect 109 -40 111 -38
rect 105 -41 111 -40
rect 149 -39 151 -37
rect 153 -39 155 -37
rect 149 -40 155 -39
rect 168 -37 174 -31
rect 168 -39 170 -37
rect 172 -39 174 -37
rect 168 -40 174 -39
rect 211 -38 217 -31
rect 255 -37 261 -31
rect 211 -40 213 -38
rect 215 -40 217 -38
rect 211 -41 217 -40
rect 255 -39 257 -37
rect 259 -39 261 -37
rect 255 -40 261 -39
rect 274 -37 280 -31
rect 274 -39 276 -37
rect 278 -39 280 -37
rect 274 -40 280 -39
rect 317 -38 323 -31
rect 361 -37 367 -31
rect 317 -40 319 -38
rect 321 -40 323 -38
rect 317 -41 323 -40
rect 361 -39 363 -37
rect 365 -39 367 -37
rect 361 -40 367 -39
rect 380 -37 386 -31
rect 380 -39 382 -37
rect 384 -39 386 -37
rect 380 -40 386 -39
rect 423 -38 429 -31
rect 467 -37 473 -31
rect 423 -40 425 -38
rect 427 -40 429 -38
rect 423 -41 429 -40
rect 467 -39 469 -37
rect 471 -39 473 -37
rect 467 -40 473 -39
rect 486 -37 492 -31
rect 486 -39 488 -37
rect 490 -39 492 -37
rect 486 -40 492 -39
rect 529 -38 535 -31
rect 573 -37 579 -31
rect 529 -40 531 -38
rect 533 -40 535 -38
rect 529 -41 535 -40
rect 573 -39 575 -37
rect 577 -39 579 -37
rect 573 -40 579 -39
rect 592 -37 598 -31
rect 592 -39 594 -37
rect 596 -39 598 -37
rect 592 -40 598 -39
rect 635 -38 641 -31
rect 679 -37 685 -31
rect 635 -40 637 -38
rect 639 -40 641 -38
rect 635 -41 641 -40
rect 679 -39 681 -37
rect 683 -39 685 -37
rect 679 -40 685 -39
rect 698 -37 704 -31
rect 698 -39 700 -37
rect 702 -39 704 -37
rect 698 -40 704 -39
rect 741 -38 747 -31
rect 785 -37 791 -31
rect 741 -40 743 -38
rect 745 -40 747 -38
rect 741 -41 747 -40
rect 785 -39 787 -37
rect 789 -39 791 -37
rect 785 -40 791 -39
rect 804 -37 810 -31
rect 804 -39 806 -37
rect 808 -39 810 -37
rect 804 -40 810 -39
rect 847 -38 853 -31
rect 891 -37 897 -31
rect 847 -40 849 -38
rect 851 -40 853 -38
rect 847 -41 853 -40
rect 891 -39 893 -37
rect 895 -39 897 -37
rect 891 -40 897 -39
rect 910 -37 916 -31
rect 910 -39 912 -37
rect 914 -39 916 -37
rect 910 -40 916 -39
rect -12 -46 5 -45
rect -12 -48 -10 -46
rect -8 -48 5 -46
rect -12 -49 5 -48
rect 9 -46 16 -45
rect 9 -48 11 -46
rect 13 -48 16 -46
rect 9 -49 16 -48
rect 1 -53 5 -49
rect 1 -57 9 -53
rect 5 -62 9 -57
rect 5 -64 6 -62
rect 8 -64 9 -62
rect 5 -69 9 -64
rect -9 -72 9 -69
rect -9 -74 -8 -72
rect -6 -73 9 -72
rect 12 -72 16 -49
rect -6 -74 -5 -73
rect -9 -76 -5 -74
rect 12 -74 13 -72
rect 15 -74 16 -72
rect 12 -76 16 -74
rect 27 -45 80 -44
rect 27 -47 76 -45
rect 78 -47 80 -45
rect 27 -48 80 -47
rect 27 -62 31 -48
rect 27 -64 28 -62
rect 30 -64 31 -62
rect 27 -66 31 -64
rect 34 -53 38 -51
rect 34 -55 35 -53
rect 37 -55 38 -53
rect 34 -76 38 -55
rect 50 -53 56 -51
rect 50 -55 53 -53
rect 55 -55 56 -53
rect 50 -57 56 -55
rect 50 -61 54 -57
rect 41 -62 54 -61
rect 41 -64 43 -62
rect 45 -64 54 -62
rect 41 -65 54 -64
rect 1 -77 7 -76
rect 1 -79 3 -77
rect 5 -79 7 -77
rect 1 -87 7 -79
rect 31 -77 38 -76
rect 50 -72 54 -65
rect 50 -74 56 -72
rect 50 -76 53 -74
rect 55 -76 56 -74
rect 31 -79 33 -77
rect 35 -79 38 -77
rect 31 -80 38 -79
rect 42 -79 46 -77
rect 50 -78 56 -76
rect 76 -72 80 -48
rect 94 -46 111 -45
rect 94 -48 96 -46
rect 98 -48 111 -46
rect 94 -49 111 -48
rect 115 -46 122 -45
rect 115 -48 117 -46
rect 119 -48 122 -46
rect 115 -49 122 -48
rect 107 -53 111 -49
rect 107 -57 115 -53
rect 111 -62 115 -57
rect 111 -64 112 -62
rect 114 -64 115 -62
rect 111 -69 115 -64
rect 75 -74 80 -72
rect 75 -76 76 -74
rect 78 -76 80 -74
rect 97 -72 115 -69
rect 97 -74 98 -72
rect 100 -73 115 -72
rect 118 -72 122 -49
rect 100 -74 101 -73
rect 97 -76 101 -74
rect 118 -74 119 -72
rect 121 -74 122 -72
rect 118 -76 122 -74
rect 133 -45 186 -44
rect 133 -47 182 -45
rect 184 -47 186 -45
rect 133 -48 186 -47
rect 133 -62 137 -48
rect 133 -64 134 -62
rect 136 -64 137 -62
rect 133 -66 137 -64
rect 140 -53 144 -51
rect 140 -55 141 -53
rect 143 -55 144 -53
rect 140 -76 144 -55
rect 156 -53 162 -51
rect 156 -55 159 -53
rect 161 -55 162 -53
rect 156 -57 162 -55
rect 156 -61 160 -57
rect 147 -62 160 -61
rect 147 -64 149 -62
rect 151 -64 160 -62
rect 147 -65 160 -64
rect 75 -78 80 -76
rect 107 -77 113 -76
rect 42 -81 43 -79
rect 45 -81 46 -79
rect 107 -79 109 -77
rect 111 -79 113 -77
rect 42 -87 46 -81
rect 63 -85 69 -84
rect 63 -87 65 -85
rect 67 -87 69 -85
rect 107 -87 113 -79
rect 137 -77 144 -76
rect 156 -72 160 -65
rect 156 -74 162 -72
rect 156 -76 159 -74
rect 161 -76 162 -74
rect 137 -79 139 -77
rect 141 -79 144 -77
rect 137 -80 144 -79
rect 148 -79 152 -77
rect 156 -78 162 -76
rect 182 -72 186 -48
rect 200 -46 217 -45
rect 200 -48 202 -46
rect 204 -48 217 -46
rect 200 -49 217 -48
rect 221 -46 228 -45
rect 221 -48 223 -46
rect 225 -48 228 -46
rect 221 -49 228 -48
rect 213 -53 217 -49
rect 213 -57 221 -53
rect 217 -62 221 -57
rect 217 -64 218 -62
rect 220 -64 221 -62
rect 217 -69 221 -64
rect 181 -74 186 -72
rect 181 -76 182 -74
rect 184 -76 186 -74
rect 203 -72 221 -69
rect 203 -74 204 -72
rect 206 -73 221 -72
rect 224 -72 228 -49
rect 206 -74 207 -73
rect 203 -76 207 -74
rect 224 -74 225 -72
rect 227 -74 228 -72
rect 224 -76 228 -74
rect 239 -45 292 -44
rect 239 -47 288 -45
rect 290 -47 292 -45
rect 239 -48 292 -47
rect 239 -62 243 -48
rect 239 -64 240 -62
rect 242 -64 243 -62
rect 239 -66 243 -64
rect 246 -53 250 -51
rect 246 -55 247 -53
rect 249 -55 250 -53
rect 246 -76 250 -55
rect 262 -53 268 -51
rect 262 -55 265 -53
rect 267 -55 268 -53
rect 262 -57 268 -55
rect 262 -61 266 -57
rect 253 -62 266 -61
rect 253 -64 255 -62
rect 257 -64 266 -62
rect 253 -65 266 -64
rect 181 -78 186 -76
rect 213 -77 219 -76
rect 148 -81 149 -79
rect 151 -81 152 -79
rect 213 -79 215 -77
rect 217 -79 219 -77
rect 148 -87 152 -81
rect 169 -85 175 -84
rect 169 -87 171 -85
rect 173 -87 175 -85
rect 213 -87 219 -79
rect 243 -77 250 -76
rect 262 -72 266 -65
rect 262 -74 268 -72
rect 262 -76 265 -74
rect 267 -76 268 -74
rect 243 -79 245 -77
rect 247 -79 250 -77
rect 243 -80 250 -79
rect 254 -79 258 -77
rect 262 -78 268 -76
rect 288 -72 292 -48
rect 306 -46 323 -45
rect 306 -48 308 -46
rect 310 -48 323 -46
rect 306 -49 323 -48
rect 327 -46 334 -45
rect 327 -48 329 -46
rect 331 -48 334 -46
rect 327 -49 334 -48
rect 319 -53 323 -49
rect 319 -57 327 -53
rect 323 -62 327 -57
rect 323 -64 324 -62
rect 326 -64 327 -62
rect 323 -69 327 -64
rect 287 -74 292 -72
rect 287 -76 288 -74
rect 290 -76 292 -74
rect 309 -72 327 -69
rect 309 -74 310 -72
rect 312 -73 327 -72
rect 330 -72 334 -49
rect 312 -74 313 -73
rect 309 -76 313 -74
rect 330 -74 331 -72
rect 333 -74 334 -72
rect 330 -76 334 -74
rect 345 -45 398 -44
rect 345 -47 394 -45
rect 396 -47 398 -45
rect 345 -48 398 -47
rect 345 -62 349 -48
rect 345 -64 346 -62
rect 348 -64 349 -62
rect 345 -66 349 -64
rect 352 -53 356 -51
rect 352 -55 353 -53
rect 355 -55 356 -53
rect 352 -76 356 -55
rect 368 -53 374 -51
rect 368 -55 371 -53
rect 373 -55 374 -53
rect 368 -57 374 -55
rect 368 -61 372 -57
rect 359 -62 372 -61
rect 359 -64 361 -62
rect 363 -64 372 -62
rect 359 -65 372 -64
rect 287 -78 292 -76
rect 319 -77 325 -76
rect 254 -81 255 -79
rect 257 -81 258 -79
rect 319 -79 321 -77
rect 323 -79 325 -77
rect 254 -87 258 -81
rect 275 -85 281 -84
rect 275 -87 277 -85
rect 279 -87 281 -85
rect 319 -87 325 -79
rect 349 -77 356 -76
rect 368 -72 372 -65
rect 368 -74 374 -72
rect 368 -76 371 -74
rect 373 -76 374 -74
rect 349 -79 351 -77
rect 353 -79 356 -77
rect 349 -80 356 -79
rect 360 -79 364 -77
rect 368 -78 374 -76
rect 394 -72 398 -48
rect 412 -46 429 -45
rect 412 -48 414 -46
rect 416 -48 429 -46
rect 412 -49 429 -48
rect 433 -46 440 -45
rect 433 -48 435 -46
rect 437 -48 440 -46
rect 433 -49 440 -48
rect 425 -53 429 -49
rect 425 -57 433 -53
rect 429 -62 433 -57
rect 429 -64 430 -62
rect 432 -64 433 -62
rect 429 -69 433 -64
rect 393 -74 398 -72
rect 393 -76 394 -74
rect 396 -76 398 -74
rect 415 -72 433 -69
rect 415 -74 416 -72
rect 418 -73 433 -72
rect 436 -72 440 -49
rect 418 -74 419 -73
rect 415 -76 419 -74
rect 436 -74 437 -72
rect 439 -74 440 -72
rect 436 -76 440 -74
rect 451 -45 504 -44
rect 451 -47 500 -45
rect 502 -47 504 -45
rect 451 -48 504 -47
rect 451 -62 455 -48
rect 451 -64 452 -62
rect 454 -64 455 -62
rect 451 -66 455 -64
rect 458 -53 462 -51
rect 458 -55 459 -53
rect 461 -55 462 -53
rect 458 -76 462 -55
rect 474 -53 480 -51
rect 474 -55 477 -53
rect 479 -55 480 -53
rect 474 -57 480 -55
rect 474 -61 478 -57
rect 465 -62 478 -61
rect 465 -64 467 -62
rect 469 -64 478 -62
rect 465 -65 478 -64
rect 393 -78 398 -76
rect 425 -77 431 -76
rect 360 -81 361 -79
rect 363 -81 364 -79
rect 425 -79 427 -77
rect 429 -79 431 -77
rect 360 -87 364 -81
rect 381 -85 387 -84
rect 381 -87 383 -85
rect 385 -87 387 -85
rect 425 -87 431 -79
rect 455 -77 462 -76
rect 474 -72 478 -65
rect 474 -74 480 -72
rect 474 -76 477 -74
rect 479 -76 480 -74
rect 455 -79 457 -77
rect 459 -79 462 -77
rect 455 -80 462 -79
rect 466 -79 470 -77
rect 474 -78 480 -76
rect 500 -72 504 -48
rect 518 -46 535 -45
rect 518 -48 520 -46
rect 522 -48 535 -46
rect 518 -49 535 -48
rect 539 -46 546 -45
rect 539 -48 541 -46
rect 543 -48 546 -46
rect 539 -49 546 -48
rect 531 -53 535 -49
rect 531 -57 539 -53
rect 535 -62 539 -57
rect 535 -64 536 -62
rect 538 -64 539 -62
rect 535 -69 539 -64
rect 499 -74 504 -72
rect 499 -76 500 -74
rect 502 -76 504 -74
rect 521 -72 539 -69
rect 521 -74 522 -72
rect 524 -73 539 -72
rect 542 -72 546 -49
rect 524 -74 525 -73
rect 521 -76 525 -74
rect 542 -74 543 -72
rect 545 -74 546 -72
rect 542 -76 546 -74
rect 557 -45 610 -44
rect 557 -47 606 -45
rect 608 -47 610 -45
rect 557 -48 610 -47
rect 557 -62 561 -48
rect 557 -64 558 -62
rect 560 -64 561 -62
rect 557 -66 561 -64
rect 564 -53 568 -51
rect 564 -55 565 -53
rect 567 -55 568 -53
rect 564 -76 568 -55
rect 580 -53 586 -51
rect 580 -55 583 -53
rect 585 -55 586 -53
rect 580 -57 586 -55
rect 580 -61 584 -57
rect 571 -62 584 -61
rect 571 -64 573 -62
rect 575 -64 584 -62
rect 571 -65 584 -64
rect 499 -78 504 -76
rect 531 -77 537 -76
rect 466 -81 467 -79
rect 469 -81 470 -79
rect 531 -79 533 -77
rect 535 -79 537 -77
rect 466 -87 470 -81
rect 487 -85 493 -84
rect 487 -87 489 -85
rect 491 -87 493 -85
rect 531 -87 537 -79
rect 561 -77 568 -76
rect 580 -72 584 -65
rect 580 -74 586 -72
rect 580 -76 583 -74
rect 585 -76 586 -74
rect 561 -79 563 -77
rect 565 -79 568 -77
rect 561 -80 568 -79
rect 572 -79 576 -77
rect 580 -78 586 -76
rect 606 -72 610 -48
rect 624 -46 641 -45
rect 624 -48 626 -46
rect 628 -48 641 -46
rect 624 -49 641 -48
rect 645 -46 652 -45
rect 645 -48 647 -46
rect 649 -48 652 -46
rect 645 -49 652 -48
rect 637 -53 641 -49
rect 637 -57 645 -53
rect 641 -62 645 -57
rect 641 -64 642 -62
rect 644 -64 645 -62
rect 641 -69 645 -64
rect 605 -74 610 -72
rect 605 -76 606 -74
rect 608 -76 610 -74
rect 627 -72 645 -69
rect 627 -74 628 -72
rect 630 -73 645 -72
rect 648 -72 652 -49
rect 630 -74 631 -73
rect 627 -76 631 -74
rect 648 -74 649 -72
rect 651 -74 652 -72
rect 648 -76 652 -74
rect 663 -45 716 -44
rect 663 -47 712 -45
rect 714 -47 716 -45
rect 663 -48 716 -47
rect 663 -62 667 -48
rect 663 -64 664 -62
rect 666 -64 667 -62
rect 663 -66 667 -64
rect 670 -53 674 -51
rect 670 -55 671 -53
rect 673 -55 674 -53
rect 670 -76 674 -55
rect 686 -53 692 -51
rect 686 -55 689 -53
rect 691 -55 692 -53
rect 686 -57 692 -55
rect 686 -61 690 -57
rect 677 -62 690 -61
rect 677 -64 679 -62
rect 681 -64 690 -62
rect 677 -65 690 -64
rect 605 -78 610 -76
rect 637 -77 643 -76
rect 572 -81 573 -79
rect 575 -81 576 -79
rect 637 -79 639 -77
rect 641 -79 643 -77
rect 572 -87 576 -81
rect 593 -85 599 -84
rect 593 -87 595 -85
rect 597 -87 599 -85
rect 637 -87 643 -79
rect 667 -77 674 -76
rect 686 -72 690 -65
rect 686 -74 692 -72
rect 686 -76 689 -74
rect 691 -76 692 -74
rect 667 -79 669 -77
rect 671 -79 674 -77
rect 667 -80 674 -79
rect 678 -79 682 -77
rect 686 -78 692 -76
rect 712 -72 716 -48
rect 730 -46 747 -45
rect 730 -48 732 -46
rect 734 -48 747 -46
rect 730 -49 747 -48
rect 751 -46 758 -45
rect 751 -48 753 -46
rect 755 -48 758 -46
rect 751 -49 758 -48
rect 743 -53 747 -49
rect 743 -57 751 -53
rect 747 -62 751 -57
rect 747 -64 748 -62
rect 750 -64 751 -62
rect 747 -69 751 -64
rect 711 -74 716 -72
rect 711 -76 712 -74
rect 714 -76 716 -74
rect 733 -72 751 -69
rect 733 -74 734 -72
rect 736 -73 751 -72
rect 754 -72 758 -49
rect 736 -74 737 -73
rect 733 -76 737 -74
rect 754 -74 755 -72
rect 757 -74 758 -72
rect 754 -76 758 -74
rect 769 -45 822 -44
rect 769 -47 818 -45
rect 820 -47 822 -45
rect 769 -48 822 -47
rect 769 -62 773 -48
rect 769 -64 770 -62
rect 772 -64 773 -62
rect 769 -66 773 -64
rect 776 -53 780 -51
rect 776 -55 777 -53
rect 779 -55 780 -53
rect 776 -76 780 -55
rect 792 -53 798 -51
rect 792 -55 795 -53
rect 797 -55 798 -53
rect 792 -57 798 -55
rect 792 -61 796 -57
rect 783 -62 796 -61
rect 783 -64 785 -62
rect 787 -64 796 -62
rect 783 -65 796 -64
rect 711 -78 716 -76
rect 743 -77 749 -76
rect 678 -81 679 -79
rect 681 -81 682 -79
rect 743 -79 745 -77
rect 747 -79 749 -77
rect 678 -87 682 -81
rect 699 -85 705 -84
rect 699 -87 701 -85
rect 703 -87 705 -85
rect 743 -87 749 -79
rect 773 -77 780 -76
rect 792 -72 796 -65
rect 792 -74 798 -72
rect 792 -76 795 -74
rect 797 -76 798 -74
rect 773 -79 775 -77
rect 777 -79 780 -77
rect 773 -80 780 -79
rect 784 -79 788 -77
rect 792 -78 798 -76
rect 818 -72 822 -48
rect 836 -46 853 -45
rect 836 -48 838 -46
rect 840 -48 853 -46
rect 836 -49 853 -48
rect 857 -46 864 -45
rect 857 -48 859 -46
rect 861 -48 864 -46
rect 857 -49 864 -48
rect 817 -74 822 -72
rect 817 -76 818 -74
rect 820 -76 822 -74
rect 817 -78 822 -76
rect 784 -81 785 -79
rect 787 -81 788 -79
rect 784 -87 788 -81
rect 805 -85 811 -84
rect 805 -87 807 -85
rect 809 -87 811 -85
rect 849 -53 853 -49
rect 849 -57 857 -53
rect 853 -62 857 -57
rect 853 -64 854 -62
rect 856 -64 857 -62
rect 853 -69 857 -64
rect 839 -72 857 -69
rect 839 -74 840 -72
rect 842 -73 857 -72
rect 860 -72 864 -49
rect 842 -74 843 -73
rect 839 -76 843 -74
rect 860 -74 861 -72
rect 863 -74 864 -72
rect 860 -76 864 -74
rect 875 -45 928 -44
rect 875 -47 924 -45
rect 926 -47 928 -45
rect 875 -48 928 -47
rect 875 -62 879 -48
rect 875 -64 876 -62
rect 878 -64 879 -62
rect 875 -66 879 -64
rect 882 -53 886 -51
rect 882 -55 883 -53
rect 885 -55 886 -53
rect 882 -76 886 -55
rect 898 -53 904 -51
rect 898 -55 901 -53
rect 903 -55 904 -53
rect 898 -57 904 -55
rect 898 -61 902 -57
rect 889 -62 902 -61
rect 889 -64 891 -62
rect 893 -64 902 -62
rect 889 -65 902 -64
rect 849 -77 855 -76
rect 849 -79 851 -77
rect 853 -79 855 -77
rect 849 -87 855 -79
rect 879 -77 886 -76
rect 898 -72 902 -65
rect 898 -74 904 -72
rect 898 -76 901 -74
rect 903 -76 904 -74
rect 879 -79 881 -77
rect 883 -79 886 -77
rect 879 -80 886 -79
rect 890 -79 894 -77
rect 898 -78 904 -76
rect 924 -72 928 -48
rect 923 -74 928 -72
rect 923 -76 924 -74
rect 926 -76 928 -74
rect 923 -78 928 -76
rect 890 -81 891 -79
rect 893 -81 894 -79
rect 890 -87 894 -81
rect 911 -85 917 -84
rect 911 -87 913 -85
rect 915 -87 917 -85
<< via1 >>
rect 89 1163 91 1165
rect 137 1164 139 1166
rect 81 1140 83 1142
rect 133 1139 135 1141
rect 193 1170 195 1172
rect 165 1164 167 1166
rect 165 1147 167 1149
rect 210 1161 212 1163
rect 237 1164 239 1166
rect 154 1134 156 1136
rect 217 1138 219 1140
rect 285 1161 287 1163
rect 235 1130 237 1132
rect 299 1172 301 1174
rect 323 1164 325 1166
rect 307 1158 309 1160
rect 339 1161 341 1163
rect 339 1146 341 1148
rect 374 1156 376 1158
rect 367 1138 369 1140
rect 591 1147 593 1149
rect 574 1139 576 1141
rect 661 1160 663 1162
rect 621 1154 623 1156
rect 605 1130 607 1132
rect 684 1164 686 1166
rect 730 1171 732 1173
rect 730 1163 732 1165
rect 707 1146 709 1148
rect 740 1147 742 1149
rect 682 1140 684 1142
rect 145 1089 147 1091
rect 105 1084 107 1086
rect 81 1068 83 1070
rect 97 1066 99 1068
rect 133 1076 135 1078
rect 117 1058 119 1060
rect 168 1083 170 1085
rect 198 1091 200 1093
rect 169 1069 171 1071
rect 257 1099 259 1101
rect 221 1083 223 1085
rect 265 1091 267 1093
rect 213 1066 215 1068
rect 230 1066 232 1068
rect 582 1091 584 1093
rect 273 1083 275 1085
rect 574 1074 576 1076
rect 298 1067 300 1069
rect 321 1068 323 1070
rect 634 1092 636 1094
rect 602 1081 604 1083
rect 655 1084 657 1086
rect 627 1066 629 1068
rect 664 1067 666 1069
rect 672 1058 674 1060
rect 691 1092 693 1094
rect 740 1091 742 1093
rect 684 1067 686 1069
rect 732 1066 734 1068
rect 89 1019 91 1021
rect 137 1018 139 1020
rect 81 996 83 998
rect 204 1027 206 1029
rect 161 1018 163 1020
rect 196 1019 198 1021
rect 168 1002 170 1004
rect 237 1003 239 1005
rect 305 1027 307 1029
rect 273 1019 275 1021
rect 290 1011 292 1013
rect 149 994 151 996
rect 245 995 247 997
rect 272 995 274 997
rect 512 1028 514 1030
rect 606 1019 608 1021
rect 528 1012 530 1014
rect 556 1011 558 1013
rect 636 1019 638 1021
rect 628 1003 630 1005
rect 598 997 600 999
rect 715 1019 717 1021
rect 688 1011 690 1013
rect 674 999 676 1001
rect 707 1002 709 1004
rect 663 995 665 997
rect 724 998 726 1000
rect 105 940 107 942
rect 105 932 107 934
rect 81 922 83 924
rect 177 947 179 949
rect 78 914 80 916
rect 125 922 127 924
rect 145 923 147 925
rect 117 914 119 916
rect 249 955 251 957
rect 201 932 203 934
rect 185 914 187 916
rect 269 948 271 950
rect 240 923 242 925
rect 300 944 302 946
rect 277 922 279 924
rect 567 956 569 958
rect 512 924 514 926
rect 612 947 614 949
rect 558 923 560 925
rect 580 923 582 925
rect 689 947 691 949
rect 644 939 646 941
rect 605 931 607 933
rect 627 931 629 933
rect 672 932 674 934
rect 740 947 742 949
rect 732 923 734 925
rect 684 915 686 917
rect 78 876 80 878
rect 106 876 108 878
rect 97 863 99 865
rect 141 876 143 878
rect 140 859 142 861
rect 117 845 119 847
rect 190 873 192 875
rect 166 854 168 856
rect 229 867 231 869
rect 198 850 200 852
rect 251 862 253 864
rect 219 851 221 853
rect 265 873 267 875
rect 281 866 283 868
rect 317 876 319 878
rect 293 854 295 856
rect 325 859 327 861
rect 378 876 380 878
rect 361 867 363 869
rect 504 867 506 869
rect 338 843 340 845
rect 370 851 372 853
rect 519 876 521 878
rect 487 850 489 852
rect 540 876 542 878
rect 567 876 569 878
rect 560 858 562 860
rect 540 850 542 852
rect 592 853 594 855
rect 609 853 611 855
rect 623 867 625 869
rect 655 871 657 873
rect 704 884 706 886
rect 681 867 683 869
rect 696 865 698 867
rect 724 875 726 877
rect 640 850 642 852
rect 664 852 666 854
rect 708 850 710 852
rect 719 847 721 849
rect 102 807 104 809
rect 113 804 115 806
rect 97 779 99 781
rect 157 802 159 804
rect 181 804 183 806
rect 140 787 142 789
rect 117 770 119 772
rect 166 783 168 785
rect 198 787 200 789
rect 212 801 214 803
rect 125 770 127 772
rect 229 801 231 803
rect 281 804 283 806
rect 261 796 263 798
rect 254 778 256 780
rect 281 778 283 780
rect 334 804 336 806
rect 302 778 304 780
rect 451 803 453 805
rect 483 811 485 813
rect 317 787 319 789
rect 460 787 462 789
rect 443 778 445 780
rect 496 795 498 797
rect 528 800 530 802
rect 504 778 506 780
rect 540 788 542 790
rect 556 781 558 783
rect 602 803 604 805
rect 570 792 572 794
rect 623 804 625 806
rect 592 787 594 789
rect 655 800 657 802
rect 631 781 633 783
rect 704 809 706 811
rect 681 795 683 797
rect 680 778 682 780
rect 724 791 726 793
rect 715 778 717 780
rect 743 778 745 780
rect 137 739 139 741
rect 89 731 91 733
rect 81 709 83 711
rect 149 722 151 724
rect 194 723 196 725
rect 216 723 218 725
rect 177 715 179 717
rect 132 707 134 709
rect 241 731 243 733
rect 263 731 265 733
rect 209 707 211 709
rect 309 729 311 731
rect 254 698 256 700
rect 329 731 331 733
rect 544 732 546 734
rect 329 707 331 709
rect 521 710 523 712
rect 581 731 583 733
rect 552 706 554 708
rect 636 740 638 742
rect 620 721 622 723
rect 572 699 574 701
rect 704 740 706 742
rect 676 731 678 733
rect 696 732 698 734
rect 743 740 745 742
rect 644 707 646 709
rect 740 732 742 734
rect 716 722 718 724
rect 716 714 718 716
rect 97 656 99 658
rect 158 659 160 661
rect 114 652 116 654
rect 147 655 149 657
rect 133 643 135 645
rect 106 635 108 637
rect 223 657 225 659
rect 193 651 195 653
rect 185 635 187 637
rect 265 643 267 645
rect 215 635 217 637
rect 549 659 551 661
rect 576 659 578 661
rect 672 660 674 662
rect 531 643 533 645
rect 548 635 550 637
rect 516 627 518 629
rect 584 651 586 653
rect 653 652 655 654
rect 625 635 627 637
rect 660 636 662 638
rect 617 627 619 629
rect 740 660 742 662
rect 684 636 686 638
rect 732 635 734 637
rect 89 588 91 590
rect 137 587 139 589
rect 81 565 83 567
rect 130 562 132 564
rect 149 596 151 598
rect 157 587 159 589
rect 194 588 196 590
rect 166 570 168 572
rect 219 573 221 575
rect 187 562 189 564
rect 500 586 502 588
rect 523 587 525 589
rect 247 580 249 582
rect 548 571 550 573
rect 239 563 241 565
rect 591 588 593 590
rect 608 588 610 590
rect 556 563 558 565
rect 600 571 602 573
rect 564 555 566 557
rect 652 585 654 587
rect 623 563 625 565
rect 653 571 655 573
rect 704 596 706 598
rect 688 578 690 580
rect 724 588 726 590
rect 740 586 742 588
rect 716 570 718 572
rect 676 565 678 567
rect 139 514 141 516
rect 81 507 83 509
rect 114 508 116 510
rect 91 491 93 493
rect 91 483 93 485
rect 137 490 139 492
rect 216 524 218 526
rect 200 500 202 502
rect 160 495 162 497
rect 247 515 249 517
rect 239 507 241 509
rect 454 516 456 518
rect 447 498 449 500
rect 482 508 484 510
rect 482 493 484 495
rect 514 496 516 498
rect 498 490 500 492
rect 522 482 524 484
rect 586 524 588 526
rect 536 493 538 495
rect 604 516 606 518
rect 667 520 669 522
rect 584 490 586 492
rect 611 493 613 495
rect 656 507 658 509
rect 656 490 658 492
rect 628 484 630 486
rect 688 515 690 517
rect 740 514 742 516
rect 684 490 686 492
rect 732 491 734 493
rect 6 333 8 335
rect 6 323 8 325
rect 78 340 80 342
rect 178 348 180 350
rect 86 339 88 341
rect 106 324 108 326
rect 138 320 140 322
rect 186 339 188 341
rect 202 347 204 349
rect 206 323 208 325
rect 238 327 240 329
rect 278 347 280 349
rect 286 339 288 341
rect 306 331 308 333
rect 307 323 309 325
rect 338 323 340 325
rect 386 339 388 341
rect 386 323 388 325
rect 406 323 408 325
rect 438 319 440 321
rect 486 339 488 341
rect 478 329 480 331
rect 501 347 503 349
rect 538 331 540 333
rect 601 348 603 350
rect 586 339 588 341
rect 586 323 588 325
rect 606 326 608 328
rect 638 331 640 333
rect 686 339 688 341
rect 686 323 688 325
rect 702 347 704 349
rect 706 323 708 325
rect 786 339 788 341
rect 786 323 788 325
rect 29 308 31 310
rect 729 308 731 310
rect 22 254 24 256
rect 14 245 16 247
rect 63 237 65 239
rect 99 237 101 239
rect 114 262 116 264
rect 114 245 116 247
rect 199 261 201 263
rect 191 254 193 256
rect 222 254 224 256
rect 214 245 216 247
rect 163 237 165 239
rect 299 262 301 264
rect 314 262 316 264
rect 314 245 316 247
rect 263 237 265 239
rect 391 254 393 256
rect 363 237 365 239
rect 401 237 403 239
rect 424 254 426 256
rect 416 245 418 247
rect 501 262 503 264
rect 516 262 518 264
rect 516 245 518 247
rect 465 237 467 239
rect 593 254 595 256
rect 624 254 626 256
rect 616 245 618 247
rect 565 237 567 239
rect 701 262 703 264
rect 716 262 718 264
rect 716 245 718 247
rect 665 237 667 239
rect 793 254 795 256
rect 765 237 767 239
rect 14 195 16 197
rect 99 203 101 205
rect 14 179 16 181
rect 114 195 116 197
rect 122 187 124 189
rect 62 169 64 171
rect 194 179 196 181
rect 214 195 216 197
rect 298 204 300 206
rect 214 179 216 181
rect 294 187 296 189
rect 314 195 316 197
rect 322 187 324 189
rect 393 206 395 208
rect 393 179 395 181
rect 416 195 418 197
rect 416 179 418 181
rect 496 187 498 189
rect 516 195 518 197
rect 524 187 526 189
rect 596 179 598 181
rect 616 195 618 197
rect 616 179 618 181
rect 696 187 698 189
rect 716 195 718 197
rect 724 187 726 189
rect 811 189 813 191
rect 795 179 797 181
rect 171 164 173 166
rect 271 164 273 166
rect 371 164 373 166
rect 473 164 475 166
rect 573 164 575 166
rect 673 164 675 166
rect 773 164 775 166
rect 14 117 16 119
rect 62 113 64 115
rect 94 117 96 119
rect 122 109 124 111
rect 23 92 25 94
rect 262 128 264 130
rect 162 101 164 103
rect 198 117 200 119
rect 122 92 124 94
rect 222 101 224 103
rect 294 117 296 119
rect 294 109 296 111
rect 314 117 316 119
rect 222 92 224 94
rect 362 109 364 111
rect 394 117 396 119
rect 416 117 418 119
rect 322 92 324 94
rect 564 128 566 130
rect 664 128 666 130
rect 464 121 466 123
rect 496 117 498 119
rect 524 110 526 112
rect 424 92 426 94
rect 600 101 602 103
rect 616 118 618 120
rect 525 92 527 94
rect 701 117 703 119
rect 693 110 695 112
rect 625 92 627 94
rect 724 104 726 106
rect 764 96 766 98
rect 795 117 797 119
rect 811 117 813 119
rect 725 92 727 94
rect 6 35 8 37
rect 78 52 80 54
rect 178 60 180 62
rect 86 51 88 53
rect 106 36 108 38
rect 138 42 140 44
rect 186 51 188 53
rect 206 35 208 37
rect 238 39 240 41
rect 278 59 280 61
rect 286 51 288 53
rect 306 43 308 45
rect 338 32 340 34
rect 386 51 388 53
rect 386 35 388 37
rect 406 35 408 37
rect 438 31 440 33
rect 486 51 488 53
rect 478 41 480 43
rect 501 59 503 61
rect 506 43 508 45
rect 538 31 540 33
rect 601 60 603 62
rect 586 51 588 53
rect 586 35 588 37
rect 638 25 640 27
rect 686 51 688 53
rect 686 35 688 37
rect 702 59 704 61
rect 738 31 740 33
rect 786 51 788 53
rect 786 35 788 37
rect 29 20 31 22
rect -11 -64 -9 -62
rect 68 -56 70 -54
rect 95 -55 97 -53
rect 174 -56 176 -54
rect 61 -80 63 -78
rect 201 -56 203 -54
rect 280 -56 282 -54
rect 167 -80 169 -78
rect 307 -55 309 -53
rect 386 -56 388 -54
rect 273 -80 275 -78
rect 413 -56 415 -54
rect 491 -57 493 -55
rect 379 -80 381 -78
rect 519 -56 521 -54
rect 598 -56 600 -54
rect 485 -80 487 -78
rect 625 -56 627 -54
rect 702 -56 704 -54
rect 591 -80 593 -78
rect 731 -57 733 -55
rect 809 -56 811 -54
rect 697 -80 699 -78
rect 803 -80 805 -78
rect 916 -56 918 -54
rect 909 -80 911 -78
<< via2 >>
rect 315 1164 317 1166
rect 81 1053 83 1055
rect 51 1011 53 1013
rect 285 1161 287 1163
rect 348 1161 350 1163
rect 210 1157 212 1159
rect 51 983 53 985
rect 81 926 83 928
rect 51 720 53 722
rect 661 1160 663 1162
rect 145 1105 147 1107
rect 164 1083 166 1085
rect 174 1069 176 1071
rect 202 1105 204 1107
rect 337 1105 339 1107
rect 213 1045 215 1047
rect 230 1069 232 1071
rect 345 1060 347 1062
rect 337 1052 339 1054
rect 221 1045 223 1047
rect 157 1035 159 1037
rect 134 1026 136 1028
rect 370 1011 372 1013
rect 149 961 151 963
rect 272 991 274 993
rect 149 947 151 949
rect 272 948 274 950
rect 309 948 311 950
rect 201 932 203 934
rect 105 922 107 924
rect 121 922 123 924
rect 270 922 272 924
rect 121 899 123 901
rect 345 899 347 901
rect 149 889 151 891
rect 325 889 327 891
rect 157 881 159 883
rect 113 837 115 839
rect 117 795 119 797
rect 32 717 34 719
rect 51 701 53 703
rect 32 690 34 692
rect 32 587 34 589
rect 21 580 23 582
rect 97 775 99 777
rect 181 881 183 883
rect 221 873 223 875
rect 255 873 257 875
rect 204 850 206 852
rect 181 837 183 839
rect 198 817 200 819
rect 270 837 272 839
rect 281 817 283 819
rect 276 796 278 798
rect 125 745 127 747
rect 263 745 265 747
rect 309 729 311 731
rect 185 621 187 623
rect 276 681 278 683
rect 247 621 249 623
rect 257 605 259 607
rect 185 596 187 598
rect 51 579 53 581
rect 21 552 23 554
rect 32 550 34 552
rect 51 551 53 553
rect 81 549 83 551
rect 247 575 249 577
rect 370 630 372 632
rect 378 621 380 623
rect 443 1033 445 1035
rect 451 1024 453 1026
rect 556 1105 558 1107
rect 574 1079 576 1081
rect 740 1105 742 1107
rect 766 1091 768 1093
rect 636 1058 638 1060
rect 564 1049 566 1051
rect 574 1033 576 1035
rect 545 973 547 975
rect 636 1033 638 1035
rect 512 924 514 926
rect 545 858 547 860
rect 540 837 542 839
rect 551 817 553 819
rect 623 837 625 839
rect 640 817 642 819
rect 617 804 619 806
rect 566 781 568 783
rect 600 781 602 783
rect 640 773 642 775
rect 696 865 698 867
rect 724 879 726 881
rect 704 859 706 861
rect 708 817 710 819
rect 664 773 666 775
rect 496 765 498 767
rect 672 765 674 767
rect 476 755 478 757
rect 700 755 702 757
rect 551 732 553 734
rect 700 732 702 734
rect 716 732 718 734
rect 620 721 622 723
rect 512 706 514 708
rect 549 706 551 708
rect 672 707 674 709
rect 549 663 551 665
rect 672 693 674 695
rect 451 643 453 645
rect 265 549 267 551
rect 687 628 689 630
rect 664 619 666 621
rect 600 609 602 611
rect 484 602 486 604
rect 476 594 478 596
rect 591 585 593 587
rect 608 609 610 611
rect 484 549 486 551
rect 619 549 621 551
rect 647 585 649 587
rect 657 571 659 573
rect 676 549 678 551
rect 160 495 162 497
rect 740 728 742 730
rect 611 497 613 499
rect 473 493 475 495
rect 536 493 538 495
rect 740 601 742 603
rect 506 490 508 492
rect 706 455 708 457
rect 630 433 632 435
rect 501 420 503 422
rect 100 376 102 378
rect 267 380 269 382
rect 202 372 204 374
rect 202 347 204 349
rect 501 347 503 349
rect 819 339 821 341
rect 100 331 102 333
rect 298 327 300 329
rect 597 331 599 333
rect 606 326 608 328
rect 29 302 31 304
rect 138 313 140 315
rect 307 323 309 325
rect 406 323 408 325
rect 438 323 440 325
rect 338 318 340 320
rect 638 326 640 328
rect 706 323 708 325
rect 729 302 731 304
rect 338 286 340 288
rect 701 286 703 288
rect 199 270 201 272
rect 299 270 301 272
rect 496 262 498 264
rect 701 270 703 272
rect 597 254 599 256
rect 787 254 789 256
rect 99 233 101 235
rect 263 220 265 222
rect 401 230 403 232
rect 501 226 503 228
rect 565 226 567 228
rect 665 218 667 220
rect 765 219 767 221
rect 401 206 403 208
rect 811 219 813 221
rect 401 187 403 189
rect 501 187 503 189
rect 700 187 702 189
rect 201 179 203 181
rect 601 179 603 181
rect 198 164 200 166
rect 298 164 300 166
rect 401 164 403 166
rect 94 154 96 156
rect 701 164 703 166
rect 573 154 575 156
rect 773 154 775 156
rect 198 138 200 140
rect 94 135 96 137
rect 262 121 264 123
rect 298 117 300 119
rect 496 138 498 140
rect 350 109 352 111
rect 504 130 506 132
rect 464 109 466 111
rect 604 130 606 132
rect 701 136 703 138
rect 664 120 666 122
rect 811 154 813 156
rect 62 100 64 102
rect 206 101 208 103
rect 6 86 8 88
rect 402 84 404 86
rect 604 84 606 86
rect 464 67 466 69
rect 819 51 821 53
rect 138 42 140 44
rect 206 43 208 45
rect 29 20 31 22
rect 302 43 304 45
rect 238 39 240 41
rect 402 35 404 37
rect 338 32 340 34
rect 438 31 440 33
rect 538 31 540 33
rect 664 35 666 37
rect 638 25 640 27
rect 738 31 740 33
rect 350 14 352 16
rect 95 -5 97 -3
rect 68 -56 70 -54
rect 174 -56 176 -54
rect 201 -56 203 -54
rect 280 -56 282 -54
rect 307 -55 309 -53
rect 386 -56 388 -54
rect 413 -56 415 -54
rect 491 -57 493 -55
rect 519 -56 521 -54
rect 598 -56 600 -54
rect 625 -56 627 -54
rect 702 -56 704 -54
rect 731 -57 733 -55
rect 809 -56 811 -54
rect 916 -56 918 -54
rect -11 -64 -9 -62
<< via3 >>
rect 285 1161 287 1163
rect 201 932 203 934
rect 661 1160 663 1162
rect 309 729 311 731
rect 512 924 514 926
rect 696 865 698 867
rect 160 495 162 497
rect 620 721 622 723
rect 536 493 538 495
rect 706 455 708 457
rect 691 445 693 447
rect 267 380 269 382
rect 307 323 309 325
rect 406 323 408 325
rect 706 323 708 325
rect 68 -114 70 -112
rect 174 -169 176 -167
rect 281 -186 283 -184
rect 387 -210 389 -208
rect 808 -188 810 -186
rect 702 -217 704 -215
rect 916 -261 918 -259
rect 598 -270 600 -268
rect 491 -280 493 -278
<< labels >>
rlabel alu1 15 261 15 261 1 a10
rlabel alu1 63 257 63 257 1 z0
rlabel alu1 95 257 95 257 1 a00
rlabel alu1 163 257 163 257 1 z4
rlabel alu1 195 257 195 257 1 a04
rlabel alu1 115 261 115 261 1 a14
rlabel alu1 215 261 215 261 1 a12
rlabel alu1 263 257 263 257 1 z2
rlabel alu1 295 257 295 257 1 a02
rlabel alu1 315 261 315 261 1 a16
rlabel alu1 363 257 363 257 1 z6
rlabel alu1 395 257 395 257 1 a06
rlabel alu1 15 181 15 181 1 b10
rlabel alu1 63 185 63 185 1 y0
rlabel alu1 95 187 95 187 1 b00
rlabel alu1 115 181 115 181 1 b12
rlabel alu1 163 185 163 185 1 y2
rlabel alu1 195 185 195 185 1 b02
rlabel alu1 215 181 215 181 1 b14
rlabel alu1 263 185 263 185 1 y4
rlabel alu1 295 185 295 185 1 b04
rlabel alu1 315 181 315 181 1 b16
rlabel alu1 363 185 363 185 1 y6
rlabel alu1 395 185 395 185 1 b06
rlabel alu1 453 225 453 225 4 vss
rlabel alu1 453 153 453 153 2 vdd
rlabel alu1 453 81 453 81 4 vss
rlabel alu1 465 257 465 257 1 z1
rlabel alu1 497 257 497 257 1 a01
rlabel alu1 565 257 565 257 1 z5
rlabel alu1 597 257 597 257 1 a05
rlabel alu1 617 261 617 261 1 a13
rlabel alu1 665 257 665 257 1 z3
rlabel alu1 697 257 697 257 1 a03
rlabel alu1 717 261 717 261 1 a17
rlabel alu1 765 257 765 257 1 z7
rlabel alu1 797 257 797 257 1 a07
rlabel alu1 517 261 517 261 1 a15
rlabel alu1 417 261 417 261 1 a11
rlabel alu1 797 185 797 185 1 b07
rlabel alu1 765 185 765 185 1 y7
rlabel alu1 717 181 717 181 1 b17
rlabel alu1 697 185 697 185 1 b05
rlabel alu1 665 185 665 185 1 y5
rlabel alu1 618 181 618 181 1 b15
rlabel alu1 597 185 597 185 1 b03
rlabel alu1 565 185 565 185 1 y3
rlabel alu1 517 181 517 181 1 b13
rlabel alu1 417 181 417 181 1 b11
rlabel alu1 465 185 465 185 1 y1
rlabel alu1 497 185 497 185 1 b01
rlabel alu1 15 117 15 117 1 c10
rlabel alu1 63 113 63 113 1 x0
rlabel alu1 95 113 95 113 1 c00
rlabel alu1 115 117 115 117 1 c12
rlabel alu1 163 113 163 113 1 x2
rlabel alu1 195 113 195 113 1 c02
rlabel alu1 215 117 215 117 1 c13
rlabel alu1 263 113 263 113 1 x3
rlabel alu1 295 113 295 113 1 c03
rlabel alu1 315 117 315 117 1 c11
rlabel alu1 363 113 363 113 1 x1
rlabel alu1 395 113 395 113 1 c01
rlabel alu1 417 117 417 117 1 c16
rlabel alu1 465 113 465 113 1 x6
rlabel alu1 497 113 497 113 1 c06
rlabel alu1 517 117 517 117 1 c14
rlabel alu1 565 113 565 113 1 x4
rlabel alu1 617 117 617 117 1 c15
rlabel alu1 665 113 665 113 1 x5
rlabel alu1 697 113 697 113 1 c05
rlabel alu1 717 117 717 117 1 c17
rlabel alu1 765 113 765 113 1 x7
rlabel alu1 797 113 797 113 1 c07
rlabel alu1 453 287 453 287 1 vdd
rlabel alu2 597 113 597 113 1 c04
rlabel alu1 351 297 351 297 8 vdd
rlabel alu1 351 9 351 9 8 vdd
rlabel alu1 351 73 351 73 8 vss
rlabel alu1 39 329 39 329 1 q0
rlabel alu1 87 325 87 325 1 p10
rlabel alu1 139 329 139 329 1 q1
rlabel alu1 187 325 187 325 1 p11
rlabel alu1 239 329 239 329 1 q2
rlabel alu1 287 325 287 325 1 p12
rlabel alu1 339 329 339 329 1 q3
rlabel alu1 379 327 379 327 1 p13
rlabel alu1 439 329 439 329 1 q4
rlabel alu1 487 325 487 325 1 p14
rlabel alu1 539 329 539 329 1 q5
rlabel alu1 580 326 580 326 1 p15
rlabel alu1 639 329 639 329 1 q6
rlabel alu1 687 327 687 327 1 p16
rlabel alu1 739 329 739 329 1 q7
rlabel alu1 779 329 779 329 1 p17
rlabel alu1 7 41 7 41 1 r00
rlabel alu1 87 37 87 37 1 r10
rlabel alu1 107 41 107 41 1 r01
rlabel alu1 187 37 187 37 1 r11
rlabel alu1 207 41 207 41 1 r02
rlabel alu1 287 37 287 37 1 r12
rlabel alu1 307 41 307 41 1 r03
rlabel alu1 379 39 379 39 1 r13
rlabel alu1 407 41 407 41 1 r04
rlabel alu1 487 37 487 37 1 r14
rlabel alu1 507 41 507 41 1 r05
rlabel alu1 580 38 580 38 1 r15
rlabel alu1 607 41 607 41 1 r06
rlabel alu1 687 39 687 39 1 r16
rlabel alu1 707 41 707 41 1 r07
rlabel alu1 779 41 779 41 1 r17
rlabel via1 87 340 87 340 1 left_right
rlabel via1 87 52 87 52 1 left_right
rlabel alu1 39 42 39 42 1 out0
rlabel alu1 139 41 139 41 1 out1
rlabel alu1 239 42 239 42 1 out2
rlabel alu1 339 41 339 41 1 out3
rlabel alu1 439 41 439 41 1 out4
rlabel alu1 539 41 539 41 1 out5
rlabel alu1 639 42 639 42 1 out6
rlabel alu1 739 41 739 41 1 out7
rlabel alu1 351 361 351 361 8 vss
rlabel alu2 401 279 401 279 1 LR
rlabel alu1 330 688 330 688 8 vdd
rlabel alu1 330 752 330 752 8 vss
rlabel alu1 126 792 126 792 1 co1
rlabel alu1 163 1151 163 1151 1 A3
rlabel alu1 83 1134 83 1134 1 B3
rlabel alu1 173 1003 173 1003 1 A2
rlabel alu1 83 988 83 988 1 B2
rlabel alu1 150 733 150 733 1 A1
rlabel alu1 82 701 82 701 1 B1
rlabel alu1 82 558 82 558 1 B0
rlabel alu1 171 572 171 572 1 A0
rlabel space 76 1044 332 1188 1 PART4
rlabel space 73 900 308 1044 1 PART3
rlabel space 73 761 395 900 1 PART5
rlabel space 73 612 319 761 1 PART2
rlabel space 73 463 263 612 1 PART1
rlabel alu4 407 393 407 393 1 metal
rlabel alu2 386 614 386 614 1 xxx
rlabel alu3 388 606 388 606 1 yyy
rlabel alu1 521 976 521 976 8 vdd
rlabel alu1 521 1040 521 1040 8 vss
rlabel alu1 740 522 740 522 5 B7
rlabel alu1 660 505 660 505 5 A7
rlabel alu1 650 653 650 653 5 A6
rlabel alu1 740 668 740 668 5 B6
rlabel alu1 741 955 741 955 5 B5
rlabel alu1 673 923 673 923 5 A5
rlabel alu1 741 1098 741 1098 5 B4
rlabel alu1 652 1084 652 1084 5 A4
rlabel space 491 468 747 612 5 PART4
rlabel space 515 612 750 756 5 PART3
rlabel space 428 756 750 895 5 PART5
rlabel space 504 895 750 1044 5 PART2
rlabel space 560 1044 750 1193 5 PART1
rlabel alu2 434 1042 434 1042 5 xxx
rlabel alu3 434 1050 434 1050 5 yyy
rlabel alu1 34 -91 34 -91 6 vss
rlabel alu1 34 -27 34 -27 6 vdd
rlabel alu1 140 -91 140 -91 6 vss
rlabel alu1 140 -27 140 -27 6 vdd
rlabel alu1 246 -91 246 -91 6 vss
rlabel alu1 246 -27 246 -27 6 vdd
rlabel alu1 352 -91 352 -91 6 vss
rlabel alu1 352 -27 352 -27 6 vdd
rlabel alu1 458 -91 458 -91 6 vss
rlabel alu1 458 -27 458 -27 6 vdd
rlabel alu1 564 -91 564 -91 6 vss
rlabel alu1 564 -27 564 -27 6 vdd
rlabel alu1 670 -91 670 -91 6 vss
rlabel alu1 670 -27 670 -27 6 vdd
rlabel alu1 776 -91 776 -91 6 vss
rlabel alu1 776 -27 776 -27 6 vdd
rlabel alu4 62 495 62 495 1 s0
rlabel alu4 20 729 20 729 1 s1
rlabel alu4 62 933 62 933 1 s2
rlabel alu4 64 1161 64 1161 1 s3
rlabel alu4 838 493 838 493 1 s7
rlabel alu4 839 722 839 722 1 s6
rlabel alu4 833 924 833 924 1 s5
rlabel alu4 794 1161 794 1161 1 s4
rlabel alu4 833 866 833 866 1 cout
rlabel alu1 882 -91 882 -91 6 vss
rlabel alu1 882 -27 882 -27 6 vdd
rlabel alu4 59 -114 59 -114 1 s0
rlabel alu4 135 -168 135 -168 1 s1
rlabel alu4 196 -185 196 -185 1 s2
rlabel alu4 349 -209 349 -209 1 s3
rlabel alu4 502 -279 502 -279 1 s4
rlabel alu4 605 -269 605 -269 1 s5
rlabel alu4 708 -216 708 -216 1 s6
rlabel alu4 817 -186 817 -186 1 s7
rlabel alu4 925 -260 925 -260 1 cout
rlabel via2 -10 -63 -10 -63 1 out0
rlabel via2 69 -55 69 -55 1 s0
rlabel via1 62 -79 62 -79 1 shift_adder
rlabel via1 96 -54 96 -54 1 out1
rlabel via2 175 -55 175 -55 1 s1
rlabel via1 168 -79 168 -79 1 shift_adder
rlabel via2 202 -55 202 -55 1 out2
rlabel via2 281 -55 281 -55 1 s2
rlabel via1 274 -79 274 -79 1 shift_adder
rlabel via2 308 -54 308 -54 1 out3
rlabel via1 380 -79 380 -79 1 shift_adder
rlabel via2 387 -55 387 -55 1 s3
rlabel via2 414 -55 414 -55 1 out4
rlabel via2 492 -56 492 -56 1 s4
rlabel via1 486 -79 486 -79 1 shift_adder
rlabel via2 520 -55 520 -55 1 out5
rlabel via1 592 -79 592 -79 1 shift_adder
rlabel via2 599 -55 599 -55 1 s5
rlabel via2 626 -55 626 -55 1 out6
rlabel via2 703 -55 703 -55 1 s6
rlabel via1 698 -79 698 -79 1 shift_adder
rlabel via2 732 -56 732 -56 1 out7
rlabel via2 810 -55 810 -55 1 s7
rlabel via1 804 -79 804 -79 1 shift_adder
rlabel via2 917 -55 917 -55 1 cout
rlabel via1 910 -79 910 -79 1 shift_adder
rlabel alu1 7 330 7 330 1 B0
rlabel alu1 107 329 107 329 1 B1
rlabel alu1 207 330 207 330 1 B2
rlabel alu4 307 329 307 329 1 B3
rlabel alu4 407 329 407 329 1 B4
rlabel alu1 507 330 507 330 1 B5
rlabel alu3 607 330 607 330 1 B6
rlabel alu4 707 330 707 330 1 B7
rlabel via3 161 496 161 496 1 s0
rlabel via3 310 730 310 730 1 s1
rlabel via3 202 933 202 933 1 s2
rlabel via3 286 1162 286 1162 1 s3
rlabel via3 537 494 537 494 1 s7
rlabel via3 621 722 621 722 1 s6
rlabel via3 697 866 697 866 1 cout
rlabel via3 513 925 513 925 1 s5
rlabel via3 662 1161 662 1161 1 s4
rlabel via1 717 246 717 246 1 sh2
rlabel via1 617 246 617 246 1 sh2
rlabel via1 517 246 517 246 1 sh2
rlabel via1 417 246 417 246 1 sh2
rlabel via1 315 246 315 246 1 sh2
rlabel via1 215 246 215 246 1 sh2
rlabel via1 115 246 115 246 1 sh2
rlabel via1 15 246 15 246 1 sh2
rlabel via1 717 196 717 196 1 sh1
rlabel via1 617 196 617 196 1 sh1
rlabel via1 517 196 517 196 1 sh1
rlabel via1 417 196 417 196 1 sh1
rlabel via1 315 196 315 196 1 sh1
rlabel via1 215 196 215 196 1 sh1
rlabel via1 115 196 115 196 1 sh1
rlabel via1 15 196 15 196 1 sh1
rlabel via1 726 93 726 93 1 sh0
rlabel via1 626 93 626 93 1 sh0
rlabel via1 526 93 526 93 1 sh0
rlabel via1 425 93 425 93 1 sh0
rlabel via1 323 93 323 93 1 sh0
rlabel via1 223 93 223 93 1 sh0
rlabel via1 123 93 123 93 1 sh0
rlabel via1 24 93 24 93 1 sh0
rlabel alu1 19 -39 19 -39 1 res0
rlabel alu1 127 -42 127 -42 1 res1
rlabel alu1 232 -39 232 -39 1 res2
rlabel alu1 340 -43 340 -43 1 res3
rlabel alu1 444 -39 444 -39 1 res4
rlabel alu1 549 -39 549 -39 1 res5
rlabel alu1 656 -39 656 -39 1 res6
rlabel alu1 761 -41 763 -38 1 res7
rlabel alu1 867 -39 867 -39 1 res8
rlabel alu1 157 473 157 473 1 vss
rlabel alu1 154 539 154 539 1 vdd
rlabel alu1 148 613 149 613 1 vss
rlabel alu1 153 685 153 685 1 vdd
rlabel alu1 149 756 149 756 1 vss
rlabel alu1 154 828 154 828 1 vdd
rlabel alu1 153 896 153 896 1 vss
rlabel alu1 153 972 153 972 1 vdd
rlabel alu1 150 1043 150 1043 1 vss
rlabel alu1 149 1118 149 1118 1 vdd
rlabel alu1 145 1184 145 1184 1 vss
rlabel alu1 666 1184 666 1184 1 vss
rlabel alu1 668 1115 668 1115 1 vdd
rlabel alu1 672 1040 672 1040 1 vss
rlabel alu1 672 970 672 970 1 vdd
rlabel alu1 673 898 673 898 1 vss
rlabel alu1 669 826 669 826 1 vdd
rlabel alu1 669 759 669 759 1 vss
rlabel alu1 668 683 668 683 1 vdd
rlabel alu1 672 611 672 611 1 vss
rlabel alu1 670 537 670 537 1 vdd
rlabel alu1 678 471 678 471 1 vss
rlabel alu1 230 506 230 506 1 X
<< end >>
