magic
tech scmos
timestamp 1554073356
<< ab >>
rect 5 285 101 365
rect 5 281 104 285
rect 5 264 101 281
rect 105 264 201 365
rect 205 265 301 365
rect 305 289 401 365
rect 405 293 501 365
rect 505 293 601 365
rect 605 293 701 365
rect 705 293 801 365
rect 407 289 503 293
rect 507 289 603 293
rect 305 285 603 289
rect 5 260 104 264
rect 105 260 204 264
rect 205 261 304 265
rect 5 5 101 260
rect 105 120 201 260
rect 105 116 204 120
rect 105 5 201 116
rect 205 5 301 261
rect 305 237 401 285
rect 407 237 503 285
rect 507 237 603 285
rect 607 265 703 293
rect 607 261 706 265
rect 607 237 703 261
rect 305 233 703 237
rect 305 5 401 233
rect 407 211 503 233
rect 507 211 603 233
rect 607 211 703 233
rect 707 211 803 293
rect 402 209 803 211
rect 407 77 503 209
rect 507 77 603 209
rect 607 77 703 209
rect 707 77 803 209
rect 808 109 822 189
rect 405 5 501 77
rect 505 5 601 77
rect 605 5 701 77
rect 705 5 801 77
<< nwell >>
rect 0 298 806 333
rect 0 253 822 298
rect 0 109 822 189
rect 0 0 806 45
<< pwell >>
rect 0 333 806 370
rect 0 189 822 253
rect 0 72 822 109
rect 0 45 806 72
<< poly >>
rect 47 361 92 363
rect 47 356 49 361
rect 16 350 18 354
rect 27 351 29 356
rect 37 351 39 356
rect 57 353 59 357
rect 47 341 49 345
rect 77 352 79 357
rect 90 349 92 361
rect 147 361 192 363
rect 147 356 149 361
rect 116 350 118 354
rect 127 351 129 356
rect 137 351 139 356
rect 16 336 18 340
rect 27 336 29 340
rect 12 334 18 336
rect 12 332 14 334
rect 16 332 18 334
rect 12 330 18 332
rect 23 334 29 336
rect 37 337 39 340
rect 37 335 51 337
rect 23 332 25 334
rect 27 332 29 334
rect 23 330 29 332
rect 45 334 51 335
rect 45 332 47 334
rect 49 332 51 334
rect 14 327 16 330
rect 25 327 27 330
rect 35 327 37 331
rect 45 330 51 332
rect 57 336 59 342
rect 77 337 79 342
rect 90 339 92 342
rect 157 353 159 357
rect 147 341 149 345
rect 177 352 179 357
rect 190 349 192 361
rect 247 361 292 363
rect 247 356 249 361
rect 216 350 218 354
rect 227 351 229 356
rect 237 351 239 356
rect 86 337 92 339
rect 57 334 66 336
rect 57 332 62 334
rect 64 332 66 334
rect 57 330 66 332
rect 76 335 82 337
rect 76 333 78 335
rect 80 333 82 335
rect 86 335 88 337
rect 90 335 92 337
rect 116 336 118 340
rect 127 336 129 340
rect 86 333 92 335
rect 76 331 82 333
rect 45 327 47 330
rect 59 327 61 330
rect 77 327 79 331
rect 14 309 16 314
rect 90 319 92 333
rect 112 334 118 336
rect 112 332 114 334
rect 116 332 118 334
rect 112 330 118 332
rect 123 334 129 336
rect 137 337 139 340
rect 137 335 151 337
rect 123 332 125 334
rect 127 332 129 334
rect 123 330 129 332
rect 145 334 151 335
rect 145 332 147 334
rect 149 332 151 334
rect 114 327 116 330
rect 125 327 127 330
rect 135 327 137 331
rect 145 330 151 332
rect 157 336 159 342
rect 177 337 179 342
rect 190 339 192 342
rect 257 353 259 357
rect 247 341 249 345
rect 277 352 279 357
rect 290 349 292 361
rect 347 361 392 363
rect 347 356 349 361
rect 316 350 318 354
rect 327 351 329 356
rect 337 351 339 356
rect 186 337 192 339
rect 157 334 166 336
rect 157 332 162 334
rect 164 332 166 334
rect 157 330 166 332
rect 176 335 182 337
rect 176 333 178 335
rect 180 333 182 335
rect 186 335 188 337
rect 190 335 192 337
rect 216 336 218 340
rect 227 336 229 340
rect 186 333 192 335
rect 176 331 182 333
rect 145 327 147 330
rect 159 327 161 330
rect 177 327 179 331
rect 77 309 79 314
rect 114 309 116 314
rect 25 300 27 305
rect 35 297 37 305
rect 45 301 47 305
rect 59 301 61 305
rect 90 297 92 309
rect 190 319 192 333
rect 212 334 218 336
rect 212 332 214 334
rect 216 332 218 334
rect 212 330 218 332
rect 223 334 229 336
rect 237 337 239 340
rect 237 335 251 337
rect 223 332 225 334
rect 227 332 229 334
rect 223 330 229 332
rect 245 334 251 335
rect 245 332 247 334
rect 249 332 251 334
rect 214 327 216 330
rect 225 327 227 330
rect 235 327 237 331
rect 245 330 251 332
rect 257 336 259 342
rect 277 337 279 342
rect 290 339 292 342
rect 357 353 359 357
rect 347 341 349 345
rect 377 352 379 357
rect 390 349 392 361
rect 447 361 492 363
rect 447 356 449 361
rect 416 350 418 354
rect 427 351 429 356
rect 437 351 439 356
rect 286 337 292 339
rect 257 334 266 336
rect 257 332 262 334
rect 264 332 266 334
rect 257 330 266 332
rect 276 335 282 337
rect 276 333 278 335
rect 280 333 282 335
rect 286 335 288 337
rect 290 335 292 337
rect 316 336 318 340
rect 327 336 329 340
rect 286 333 292 335
rect 276 331 282 333
rect 245 327 247 330
rect 259 327 261 330
rect 277 327 279 331
rect 177 309 179 314
rect 214 309 216 314
rect 35 295 92 297
rect 125 300 127 305
rect 135 297 137 305
rect 145 301 147 305
rect 159 301 161 305
rect 190 297 192 309
rect 290 319 292 333
rect 312 334 318 336
rect 312 332 314 334
rect 316 332 318 334
rect 312 330 318 332
rect 323 334 329 336
rect 337 337 339 340
rect 337 335 351 337
rect 323 332 325 334
rect 327 332 329 334
rect 323 330 329 332
rect 345 334 351 335
rect 345 332 347 334
rect 349 332 351 334
rect 314 327 316 330
rect 325 327 327 330
rect 335 327 337 331
rect 345 330 351 332
rect 357 336 359 342
rect 377 337 379 342
rect 390 339 392 342
rect 457 353 459 357
rect 447 341 449 345
rect 477 352 479 357
rect 490 349 492 361
rect 547 361 592 363
rect 547 356 549 361
rect 516 350 518 354
rect 527 351 529 356
rect 537 351 539 356
rect 386 337 392 339
rect 357 334 366 336
rect 357 332 362 334
rect 364 332 366 334
rect 357 330 366 332
rect 376 335 382 337
rect 376 333 378 335
rect 380 333 382 335
rect 386 335 388 337
rect 390 335 392 337
rect 416 336 418 340
rect 427 336 429 340
rect 386 333 392 335
rect 376 331 382 333
rect 345 327 347 330
rect 359 327 361 330
rect 377 327 379 331
rect 277 309 279 314
rect 314 309 316 314
rect 135 295 192 297
rect 225 300 227 305
rect 235 297 237 305
rect 245 301 247 305
rect 259 301 261 305
rect 290 297 292 309
rect 390 319 392 333
rect 412 334 418 336
rect 412 332 414 334
rect 416 332 418 334
rect 412 330 418 332
rect 423 334 429 336
rect 437 337 439 340
rect 437 335 451 337
rect 423 332 425 334
rect 427 332 429 334
rect 423 330 429 332
rect 445 334 451 335
rect 445 332 447 334
rect 449 332 451 334
rect 414 327 416 330
rect 425 327 427 330
rect 435 327 437 331
rect 445 330 451 332
rect 457 336 459 342
rect 477 337 479 342
rect 490 339 492 342
rect 557 353 559 357
rect 547 341 549 345
rect 577 352 579 357
rect 590 349 592 361
rect 647 361 692 363
rect 647 356 649 361
rect 616 350 618 354
rect 627 351 629 356
rect 637 351 639 356
rect 486 337 492 339
rect 457 334 466 336
rect 457 332 462 334
rect 464 332 466 334
rect 457 330 466 332
rect 476 335 482 337
rect 476 333 478 335
rect 480 333 482 335
rect 486 335 488 337
rect 490 335 492 337
rect 516 336 518 340
rect 527 336 529 340
rect 486 333 492 335
rect 476 331 482 333
rect 445 327 447 330
rect 459 327 461 330
rect 477 327 479 331
rect 377 309 379 314
rect 414 309 416 314
rect 235 295 292 297
rect 325 300 327 305
rect 335 297 337 305
rect 345 301 347 305
rect 359 301 361 305
rect 390 297 392 309
rect 490 319 492 333
rect 512 334 518 336
rect 512 332 514 334
rect 516 332 518 334
rect 512 330 518 332
rect 523 334 529 336
rect 537 337 539 340
rect 537 335 551 337
rect 523 332 525 334
rect 527 332 529 334
rect 523 330 529 332
rect 545 334 551 335
rect 545 332 547 334
rect 549 332 551 334
rect 514 327 516 330
rect 525 327 527 330
rect 535 327 537 331
rect 545 330 551 332
rect 557 336 559 342
rect 577 337 579 342
rect 590 339 592 342
rect 657 353 659 357
rect 647 341 649 345
rect 677 352 679 357
rect 690 349 692 361
rect 747 361 792 363
rect 747 356 749 361
rect 716 350 718 354
rect 727 351 729 356
rect 737 351 739 356
rect 586 337 592 339
rect 557 334 566 336
rect 557 332 562 334
rect 564 332 566 334
rect 557 330 566 332
rect 576 335 582 337
rect 576 333 578 335
rect 580 333 582 335
rect 586 335 588 337
rect 590 335 592 337
rect 616 336 618 340
rect 627 336 629 340
rect 586 333 592 335
rect 576 331 582 333
rect 545 327 547 330
rect 559 327 561 330
rect 577 327 579 331
rect 477 309 479 314
rect 514 309 516 314
rect 335 295 392 297
rect 425 300 427 305
rect 435 297 437 305
rect 445 301 447 305
rect 459 301 461 305
rect 490 297 492 309
rect 590 319 592 333
rect 612 334 618 336
rect 612 332 614 334
rect 616 332 618 334
rect 612 330 618 332
rect 623 334 629 336
rect 637 337 639 340
rect 637 335 651 337
rect 623 332 625 334
rect 627 332 629 334
rect 623 330 629 332
rect 645 334 651 335
rect 645 332 647 334
rect 649 332 651 334
rect 614 327 616 330
rect 625 327 627 330
rect 635 327 637 331
rect 645 330 651 332
rect 657 336 659 342
rect 677 337 679 342
rect 690 339 692 342
rect 757 353 759 357
rect 747 341 749 345
rect 777 352 779 357
rect 790 349 792 361
rect 686 337 692 339
rect 657 334 666 336
rect 657 332 662 334
rect 664 332 666 334
rect 657 330 666 332
rect 676 335 682 337
rect 676 333 678 335
rect 680 333 682 335
rect 686 335 688 337
rect 690 335 692 337
rect 716 336 718 340
rect 727 336 729 340
rect 686 333 692 335
rect 676 331 682 333
rect 645 327 647 330
rect 659 327 661 330
rect 677 327 679 331
rect 577 309 579 314
rect 614 309 616 314
rect 435 295 492 297
rect 525 300 527 305
rect 535 297 537 305
rect 545 301 547 305
rect 559 301 561 305
rect 590 297 592 309
rect 690 319 692 333
rect 712 334 718 336
rect 712 332 714 334
rect 716 332 718 334
rect 712 330 718 332
rect 723 334 729 336
rect 737 337 739 340
rect 737 335 751 337
rect 723 332 725 334
rect 727 332 729 334
rect 723 330 729 332
rect 745 334 751 335
rect 745 332 747 334
rect 749 332 751 334
rect 714 327 716 330
rect 725 327 727 330
rect 735 327 737 331
rect 745 330 751 332
rect 757 336 759 342
rect 777 337 779 342
rect 790 339 792 342
rect 786 337 792 339
rect 757 334 766 336
rect 757 332 762 334
rect 764 332 766 334
rect 757 330 766 332
rect 776 335 782 337
rect 776 333 778 335
rect 780 333 782 335
rect 786 335 788 337
rect 790 335 792 337
rect 786 333 792 335
rect 776 331 782 333
rect 745 327 747 330
rect 759 327 761 330
rect 777 327 779 331
rect 677 309 679 314
rect 714 309 716 314
rect 535 295 592 297
rect 625 300 627 305
rect 635 297 637 305
rect 645 301 647 305
rect 659 301 661 305
rect 690 297 692 309
rect 790 319 792 333
rect 777 309 779 314
rect 635 295 692 297
rect 725 300 727 305
rect 735 297 737 305
rect 745 301 747 305
rect 759 301 761 305
rect 790 297 792 309
rect 735 295 792 297
rect 14 289 71 291
rect 14 277 16 289
rect 45 281 47 285
rect 59 281 61 285
rect 69 281 71 289
rect 79 281 81 286
rect 114 289 171 291
rect 27 272 29 277
rect 14 253 16 267
rect 114 277 116 289
rect 145 281 147 285
rect 159 281 161 285
rect 169 281 171 289
rect 179 281 181 286
rect 214 289 271 291
rect 90 272 92 277
rect 127 272 129 277
rect 27 255 29 259
rect 45 256 47 259
rect 59 256 61 259
rect 24 253 30 255
rect 14 251 20 253
rect 14 249 16 251
rect 18 249 20 251
rect 24 251 26 253
rect 28 251 30 253
rect 24 249 30 251
rect 40 254 49 256
rect 40 252 42 254
rect 44 252 49 254
rect 40 250 49 252
rect 14 247 20 249
rect 14 244 16 247
rect 27 244 29 249
rect 47 244 49 250
rect 55 254 61 256
rect 69 255 71 259
rect 79 256 81 259
rect 90 256 92 259
rect 55 252 57 254
rect 59 252 61 254
rect 55 251 61 252
rect 77 254 83 256
rect 77 252 79 254
rect 81 252 83 254
rect 55 249 69 251
rect 67 246 69 249
rect 77 250 83 252
rect 88 254 94 256
rect 88 252 90 254
rect 92 252 94 254
rect 88 250 94 252
rect 114 253 116 267
rect 214 277 216 289
rect 245 281 247 285
rect 259 281 261 285
rect 269 281 271 289
rect 279 281 281 286
rect 314 289 371 291
rect 190 272 192 277
rect 227 272 229 277
rect 127 255 129 259
rect 145 256 147 259
rect 159 256 161 259
rect 124 253 130 255
rect 114 251 120 253
rect 77 246 79 250
rect 88 246 90 250
rect 114 249 116 251
rect 118 249 120 251
rect 124 251 126 253
rect 128 251 130 253
rect 124 249 130 251
rect 140 254 149 256
rect 140 252 142 254
rect 144 252 149 254
rect 140 250 149 252
rect 114 247 120 249
rect 14 225 16 237
rect 27 229 29 234
rect 57 241 59 245
rect 47 229 49 233
rect 114 244 116 247
rect 127 244 129 249
rect 147 244 149 250
rect 155 254 161 256
rect 169 255 171 259
rect 179 256 181 259
rect 190 256 192 259
rect 155 252 157 254
rect 159 252 161 254
rect 155 251 161 252
rect 177 254 183 256
rect 177 252 179 254
rect 181 252 183 254
rect 155 249 169 251
rect 167 246 169 249
rect 177 250 183 252
rect 188 254 194 256
rect 188 252 190 254
rect 192 252 194 254
rect 188 250 194 252
rect 214 253 216 267
rect 314 277 316 289
rect 345 281 347 285
rect 359 281 361 285
rect 369 281 371 289
rect 379 281 381 286
rect 416 289 473 291
rect 290 273 292 277
rect 327 272 329 277
rect 227 255 229 259
rect 245 256 247 259
rect 259 256 261 259
rect 224 253 230 255
rect 214 251 220 253
rect 177 246 179 250
rect 188 246 190 250
rect 214 249 216 251
rect 218 249 220 251
rect 224 251 226 253
rect 228 251 230 253
rect 224 249 230 251
rect 240 254 249 256
rect 240 252 242 254
rect 244 252 249 254
rect 240 250 249 252
rect 214 247 220 249
rect 67 230 69 235
rect 77 230 79 235
rect 88 232 90 236
rect 57 225 59 230
rect 14 223 59 225
rect 114 225 116 237
rect 127 229 129 234
rect 157 241 159 245
rect 147 229 149 233
rect 214 244 216 247
rect 227 244 229 249
rect 247 244 249 250
rect 255 254 261 256
rect 269 255 271 259
rect 279 256 281 259
rect 290 256 292 259
rect 255 252 257 254
rect 259 252 261 254
rect 255 251 261 252
rect 277 254 283 256
rect 277 252 279 254
rect 281 252 283 254
rect 255 249 269 251
rect 267 246 269 249
rect 277 250 283 252
rect 288 254 294 256
rect 288 252 290 254
rect 292 252 294 254
rect 288 250 294 252
rect 314 253 316 267
rect 416 277 418 289
rect 447 281 449 285
rect 461 281 463 285
rect 471 281 473 289
rect 481 281 483 286
rect 516 289 573 291
rect 390 272 392 277
rect 429 272 431 277
rect 327 255 329 259
rect 345 256 347 259
rect 359 256 361 259
rect 324 253 330 255
rect 314 251 320 253
rect 277 246 279 250
rect 288 246 290 250
rect 314 249 316 251
rect 318 249 320 251
rect 324 251 326 253
rect 328 251 330 253
rect 324 249 330 251
rect 340 254 349 256
rect 340 252 342 254
rect 344 252 349 254
rect 340 250 349 252
rect 314 247 320 249
rect 167 230 169 235
rect 177 230 179 235
rect 188 232 190 236
rect 157 225 159 230
rect 114 223 159 225
rect 214 225 216 237
rect 227 229 229 234
rect 257 241 259 245
rect 247 229 249 233
rect 314 244 316 247
rect 327 244 329 249
rect 347 244 349 250
rect 355 254 361 256
rect 369 255 371 259
rect 379 256 381 259
rect 390 256 392 259
rect 355 252 357 254
rect 359 252 361 254
rect 355 251 361 252
rect 377 254 383 256
rect 377 252 379 254
rect 381 252 383 254
rect 355 249 369 251
rect 367 246 369 249
rect 377 250 383 252
rect 388 254 394 256
rect 388 252 390 254
rect 392 252 394 254
rect 388 250 394 252
rect 416 253 418 267
rect 516 277 518 289
rect 547 281 549 285
rect 561 281 563 285
rect 571 281 573 289
rect 581 281 583 286
rect 616 289 673 291
rect 492 273 494 277
rect 529 272 531 277
rect 429 255 431 259
rect 447 256 449 259
rect 461 256 463 259
rect 426 253 432 255
rect 416 251 422 253
rect 377 246 379 250
rect 388 246 390 250
rect 416 249 418 251
rect 420 249 422 251
rect 426 251 428 253
rect 430 251 432 253
rect 426 249 432 251
rect 442 254 451 256
rect 442 252 444 254
rect 446 252 451 254
rect 442 250 451 252
rect 416 247 422 249
rect 267 230 269 235
rect 277 230 279 235
rect 288 232 290 236
rect 257 225 259 230
rect 214 223 259 225
rect 314 225 316 237
rect 327 229 329 234
rect 357 241 359 245
rect 347 229 349 233
rect 416 244 418 247
rect 429 244 431 249
rect 449 244 451 250
rect 457 254 463 256
rect 471 255 473 259
rect 481 256 483 259
rect 492 256 494 260
rect 457 252 459 254
rect 461 252 463 254
rect 457 251 463 252
rect 479 254 485 256
rect 479 252 481 254
rect 483 252 485 254
rect 457 249 471 251
rect 469 246 471 249
rect 479 250 485 252
rect 490 254 496 256
rect 490 252 492 254
rect 494 252 496 254
rect 490 250 496 252
rect 516 253 518 267
rect 616 277 618 289
rect 647 281 649 285
rect 661 281 663 285
rect 671 281 673 289
rect 681 281 683 286
rect 716 289 773 291
rect 592 272 594 277
rect 629 272 631 277
rect 529 255 531 259
rect 547 256 549 259
rect 561 256 563 259
rect 526 253 532 255
rect 516 251 522 253
rect 479 246 481 250
rect 490 246 492 250
rect 516 249 518 251
rect 520 249 522 251
rect 526 251 528 253
rect 530 251 532 253
rect 526 249 532 251
rect 542 254 551 256
rect 542 252 544 254
rect 546 252 551 254
rect 542 250 551 252
rect 516 247 522 249
rect 367 230 369 235
rect 377 230 379 235
rect 388 232 390 236
rect 357 225 359 230
rect 314 223 359 225
rect 416 225 418 237
rect 429 229 431 234
rect 459 241 461 245
rect 449 229 451 233
rect 516 244 518 247
rect 529 244 531 249
rect 549 244 551 250
rect 557 254 563 256
rect 571 255 573 259
rect 581 256 583 259
rect 592 256 594 259
rect 557 252 559 254
rect 561 252 563 254
rect 557 251 563 252
rect 579 254 585 256
rect 579 252 581 254
rect 583 252 585 254
rect 557 249 571 251
rect 569 246 571 249
rect 579 250 585 252
rect 590 254 596 256
rect 590 252 592 254
rect 594 252 596 254
rect 590 250 596 252
rect 616 253 618 267
rect 716 277 718 289
rect 747 281 749 285
rect 761 281 763 285
rect 771 281 773 289
rect 781 281 783 286
rect 692 273 694 277
rect 729 272 731 277
rect 629 255 631 259
rect 647 256 649 259
rect 661 256 663 259
rect 626 253 632 255
rect 616 251 622 253
rect 579 246 581 250
rect 590 246 592 250
rect 616 249 618 251
rect 620 249 622 251
rect 626 251 628 253
rect 630 251 632 253
rect 626 249 632 251
rect 642 254 651 256
rect 642 252 644 254
rect 646 252 651 254
rect 642 250 651 252
rect 616 247 622 249
rect 469 230 471 235
rect 479 230 481 235
rect 490 232 492 236
rect 459 225 461 230
rect 416 223 461 225
rect 516 225 518 237
rect 529 229 531 234
rect 559 241 561 245
rect 549 229 551 233
rect 616 244 618 247
rect 629 244 631 249
rect 649 244 651 250
rect 657 254 663 256
rect 671 255 673 259
rect 681 256 683 259
rect 692 256 694 260
rect 657 252 659 254
rect 661 252 663 254
rect 657 251 663 252
rect 679 254 685 256
rect 679 252 681 254
rect 683 252 685 254
rect 657 249 671 251
rect 669 246 671 249
rect 679 250 685 252
rect 690 254 696 256
rect 690 252 692 254
rect 694 252 696 254
rect 690 250 696 252
rect 716 253 718 267
rect 792 272 794 277
rect 729 255 731 259
rect 747 256 749 259
rect 761 256 763 259
rect 726 253 732 255
rect 716 251 722 253
rect 679 246 681 250
rect 690 246 692 250
rect 716 249 718 251
rect 720 249 722 251
rect 726 251 728 253
rect 730 251 732 253
rect 726 249 732 251
rect 742 254 751 256
rect 742 252 744 254
rect 746 252 751 254
rect 742 250 751 252
rect 716 247 722 249
rect 569 230 571 235
rect 579 230 581 235
rect 590 232 592 236
rect 559 225 561 230
rect 516 223 561 225
rect 616 225 618 237
rect 629 229 631 234
rect 659 241 661 245
rect 649 229 651 233
rect 716 244 718 247
rect 729 244 731 249
rect 749 244 751 250
rect 757 254 763 256
rect 771 255 773 259
rect 781 256 783 259
rect 792 256 794 259
rect 757 252 759 254
rect 761 252 763 254
rect 757 251 763 252
rect 779 254 785 256
rect 779 252 781 254
rect 783 252 785 254
rect 757 249 771 251
rect 769 246 771 249
rect 779 250 785 252
rect 790 254 796 256
rect 790 252 792 254
rect 794 252 796 254
rect 790 250 796 252
rect 779 246 781 250
rect 790 246 792 250
rect 669 230 671 235
rect 679 230 681 235
rect 690 232 692 236
rect 659 225 661 230
rect 616 223 661 225
rect 716 225 718 237
rect 729 229 731 234
rect 759 241 761 245
rect 749 229 751 233
rect 769 230 771 235
rect 779 230 781 235
rect 790 232 792 236
rect 759 225 761 230
rect 716 223 761 225
rect 14 217 59 219
rect 14 205 16 217
rect 27 208 29 213
rect 47 209 49 213
rect 57 212 59 217
rect 114 217 159 219
rect 67 207 69 212
rect 77 207 79 212
rect 14 195 16 198
rect 14 193 20 195
rect 27 193 29 198
rect 14 191 16 193
rect 18 191 20 193
rect 14 189 20 191
rect 24 191 30 193
rect 47 192 49 198
rect 57 197 59 201
rect 88 206 90 210
rect 114 205 116 217
rect 127 208 129 213
rect 147 209 149 213
rect 157 212 159 217
rect 214 217 259 219
rect 167 207 169 212
rect 177 207 179 212
rect 67 193 69 196
rect 24 189 26 191
rect 28 189 30 191
rect 14 175 16 189
rect 24 187 30 189
rect 40 190 49 192
rect 40 188 42 190
rect 44 188 49 190
rect 27 183 29 187
rect 40 186 49 188
rect 55 191 69 193
rect 77 192 79 196
rect 88 192 90 196
rect 114 195 116 198
rect 114 193 120 195
rect 127 194 129 198
rect 55 190 61 191
rect 55 188 57 190
rect 59 188 61 190
rect 55 186 61 188
rect 77 190 83 192
rect 77 188 79 190
rect 81 188 83 190
rect 45 183 47 186
rect 59 183 61 186
rect 69 183 71 187
rect 77 186 83 188
rect 88 190 94 192
rect 88 188 90 190
rect 92 188 94 190
rect 88 186 94 188
rect 114 191 116 193
rect 118 191 120 193
rect 114 189 120 191
rect 124 192 130 194
rect 147 192 149 198
rect 157 197 159 201
rect 188 206 190 210
rect 214 205 216 217
rect 227 208 229 213
rect 247 209 249 213
rect 257 212 259 217
rect 314 217 359 219
rect 267 207 269 212
rect 277 207 279 212
rect 167 193 169 196
rect 124 190 126 192
rect 128 190 130 192
rect 79 183 81 186
rect 90 183 92 186
rect 27 165 29 170
rect 14 153 16 165
rect 114 175 116 189
rect 124 188 130 190
rect 140 190 149 192
rect 140 188 142 190
rect 144 188 149 190
rect 127 183 129 188
rect 140 186 149 188
rect 155 191 169 193
rect 177 192 179 196
rect 188 192 190 196
rect 214 195 216 198
rect 214 193 220 195
rect 227 193 229 198
rect 155 190 161 191
rect 155 188 157 190
rect 159 188 161 190
rect 155 186 161 188
rect 177 190 183 192
rect 177 188 179 190
rect 181 188 183 190
rect 145 183 147 186
rect 159 183 161 186
rect 169 183 171 187
rect 177 186 183 188
rect 188 190 194 192
rect 188 188 190 190
rect 192 188 194 190
rect 188 186 194 188
rect 214 191 216 193
rect 218 191 220 193
rect 214 189 220 191
rect 224 191 230 193
rect 247 192 249 198
rect 257 197 259 201
rect 288 206 290 210
rect 314 205 316 217
rect 327 208 329 213
rect 347 209 349 213
rect 357 212 359 217
rect 416 217 461 219
rect 367 207 369 212
rect 377 207 379 212
rect 267 193 269 196
rect 224 189 226 191
rect 228 189 230 191
rect 179 183 181 186
rect 190 183 192 186
rect 90 165 92 170
rect 127 165 129 170
rect 45 157 47 161
rect 59 157 61 161
rect 69 153 71 161
rect 79 156 81 161
rect 14 151 71 153
rect 114 153 116 165
rect 214 175 216 189
rect 224 187 230 189
rect 240 190 249 192
rect 240 188 242 190
rect 244 188 249 190
rect 227 183 229 187
rect 240 186 249 188
rect 255 191 269 193
rect 277 192 279 196
rect 288 192 290 196
rect 314 195 316 198
rect 314 193 320 195
rect 327 194 329 198
rect 255 190 261 191
rect 255 188 257 190
rect 259 188 261 190
rect 255 186 261 188
rect 277 190 283 192
rect 277 188 279 190
rect 281 188 283 190
rect 245 183 247 186
rect 259 183 261 186
rect 269 183 271 187
rect 277 186 283 188
rect 288 190 294 192
rect 288 188 290 190
rect 292 188 294 190
rect 288 186 294 188
rect 314 191 316 193
rect 318 191 320 193
rect 314 189 320 191
rect 324 192 330 194
rect 347 192 349 198
rect 357 197 359 201
rect 388 206 390 210
rect 416 205 418 217
rect 429 208 431 213
rect 449 209 451 213
rect 459 212 461 217
rect 516 217 561 219
rect 469 207 471 212
rect 479 207 481 212
rect 367 193 369 196
rect 324 190 326 192
rect 328 190 330 192
rect 279 183 281 186
rect 290 183 292 186
rect 190 165 192 170
rect 227 165 229 170
rect 145 157 147 161
rect 159 157 161 161
rect 169 153 171 161
rect 179 156 181 161
rect 114 151 171 153
rect 214 153 216 165
rect 314 175 316 189
rect 324 188 330 190
rect 340 190 349 192
rect 340 188 342 190
rect 344 188 349 190
rect 327 183 329 188
rect 340 186 349 188
rect 355 191 369 193
rect 377 192 379 196
rect 388 192 390 196
rect 416 195 418 198
rect 416 193 422 195
rect 429 193 431 198
rect 355 190 361 191
rect 355 188 357 190
rect 359 188 361 190
rect 355 186 361 188
rect 377 190 383 192
rect 377 188 379 190
rect 381 188 383 190
rect 345 183 347 186
rect 359 183 361 186
rect 369 183 371 187
rect 377 186 383 188
rect 387 190 394 192
rect 387 188 389 190
rect 391 188 394 190
rect 387 186 394 188
rect 416 191 418 193
rect 420 191 422 193
rect 416 189 422 191
rect 426 191 432 193
rect 449 192 451 198
rect 459 197 461 201
rect 490 206 492 210
rect 516 205 518 217
rect 529 208 531 213
rect 549 209 551 213
rect 559 212 561 217
rect 616 217 661 219
rect 569 207 571 212
rect 579 207 581 212
rect 469 193 471 196
rect 426 189 428 191
rect 430 189 432 191
rect 379 183 381 186
rect 390 183 392 186
rect 290 165 292 170
rect 327 165 329 170
rect 245 157 247 161
rect 259 157 261 161
rect 269 153 271 161
rect 279 156 281 161
rect 214 151 271 153
rect 314 153 316 165
rect 416 175 418 189
rect 426 187 432 189
rect 442 190 451 192
rect 442 188 444 190
rect 446 188 451 190
rect 429 183 431 187
rect 442 186 451 188
rect 457 191 471 193
rect 479 192 481 196
rect 490 192 492 196
rect 516 195 518 198
rect 516 193 522 195
rect 529 194 531 198
rect 457 190 463 191
rect 457 188 459 190
rect 461 188 463 190
rect 457 186 463 188
rect 479 190 485 192
rect 479 188 481 190
rect 483 188 485 190
rect 447 183 449 186
rect 461 183 463 186
rect 471 183 473 187
rect 479 186 485 188
rect 490 190 496 192
rect 490 188 492 190
rect 494 188 496 190
rect 490 186 496 188
rect 516 191 518 193
rect 520 191 522 193
rect 516 189 522 191
rect 526 192 532 194
rect 549 192 551 198
rect 559 197 561 201
rect 590 206 592 210
rect 616 205 618 217
rect 629 208 631 213
rect 649 209 651 213
rect 659 212 661 217
rect 716 217 761 219
rect 669 207 671 212
rect 679 207 681 212
rect 569 193 571 196
rect 526 190 528 192
rect 530 190 532 192
rect 481 183 483 186
rect 492 183 494 186
rect 390 165 392 170
rect 429 165 431 170
rect 345 157 347 161
rect 359 157 361 161
rect 369 153 371 161
rect 379 156 381 161
rect 314 151 371 153
rect 416 153 418 165
rect 516 175 518 189
rect 526 188 532 190
rect 542 190 551 192
rect 542 188 544 190
rect 546 188 551 190
rect 529 183 531 188
rect 542 186 551 188
rect 557 191 571 193
rect 579 192 581 196
rect 590 192 592 196
rect 616 195 618 198
rect 616 193 622 195
rect 629 193 631 198
rect 557 190 563 191
rect 557 188 559 190
rect 561 188 563 190
rect 557 186 563 188
rect 579 190 585 192
rect 579 188 581 190
rect 583 188 585 190
rect 547 183 549 186
rect 561 183 563 186
rect 571 183 573 187
rect 579 186 585 188
rect 590 190 596 192
rect 590 188 592 190
rect 594 188 596 190
rect 590 186 596 188
rect 616 191 618 193
rect 620 191 622 193
rect 616 189 622 191
rect 626 191 632 193
rect 649 192 651 198
rect 659 197 661 201
rect 690 206 692 210
rect 716 205 718 217
rect 729 208 731 213
rect 749 209 751 213
rect 759 212 761 217
rect 769 207 771 212
rect 779 207 781 212
rect 669 193 671 196
rect 626 189 628 191
rect 630 189 632 191
rect 581 183 583 186
rect 592 183 594 186
rect 492 165 494 170
rect 529 165 531 170
rect 447 157 449 161
rect 461 157 463 161
rect 471 153 473 161
rect 481 156 483 161
rect 416 151 473 153
rect 516 153 518 165
rect 616 175 618 189
rect 626 187 632 189
rect 642 190 651 192
rect 642 188 644 190
rect 646 188 651 190
rect 629 183 631 187
rect 642 186 651 188
rect 657 191 671 193
rect 679 192 681 196
rect 690 192 692 196
rect 716 195 718 198
rect 716 193 722 195
rect 729 194 731 198
rect 657 190 663 191
rect 657 188 659 190
rect 661 188 663 190
rect 657 186 663 188
rect 679 190 685 192
rect 679 188 681 190
rect 683 188 685 190
rect 647 183 649 186
rect 661 183 663 186
rect 671 183 673 187
rect 679 186 685 188
rect 690 190 696 192
rect 690 188 692 190
rect 694 188 696 190
rect 690 186 696 188
rect 716 191 718 193
rect 720 191 722 193
rect 716 189 722 191
rect 726 192 732 194
rect 749 192 751 198
rect 759 197 761 201
rect 790 206 792 210
rect 769 193 771 196
rect 726 190 728 192
rect 730 190 732 192
rect 681 183 683 186
rect 692 183 694 186
rect 592 165 594 170
rect 629 165 631 170
rect 547 157 549 161
rect 561 157 563 161
rect 571 153 573 161
rect 581 156 583 161
rect 516 151 573 153
rect 616 153 618 165
rect 716 175 718 189
rect 726 188 732 190
rect 742 190 751 192
rect 742 188 744 190
rect 746 188 751 190
rect 729 183 731 188
rect 742 186 751 188
rect 757 191 771 193
rect 779 192 781 196
rect 790 192 792 196
rect 757 190 763 191
rect 757 188 759 190
rect 761 188 763 190
rect 757 186 763 188
rect 779 190 785 192
rect 779 188 781 190
rect 783 188 785 190
rect 747 183 749 186
rect 761 183 763 186
rect 771 183 773 187
rect 779 186 785 188
rect 790 190 796 192
rect 790 188 792 190
rect 794 188 796 190
rect 790 186 796 188
rect 781 183 783 186
rect 792 183 794 186
rect 692 165 694 170
rect 729 165 731 170
rect 647 157 649 161
rect 661 157 663 161
rect 671 153 673 161
rect 681 156 683 161
rect 616 151 673 153
rect 716 153 718 165
rect 792 165 794 170
rect 747 157 749 161
rect 761 157 763 161
rect 771 153 773 161
rect 781 156 783 161
rect 716 151 773 153
rect 14 145 71 147
rect 14 133 16 145
rect 45 137 47 141
rect 59 137 61 141
rect 69 137 71 145
rect 79 137 81 142
rect 114 145 171 147
rect 27 128 29 133
rect 14 109 16 123
rect 114 133 116 145
rect 145 137 147 141
rect 159 137 161 141
rect 169 137 171 145
rect 179 137 181 142
rect 214 145 271 147
rect 90 128 92 133
rect 127 128 129 133
rect 27 111 29 115
rect 45 112 47 115
rect 59 112 61 115
rect 24 109 30 111
rect 14 107 20 109
rect 14 105 16 107
rect 18 105 20 107
rect 24 107 26 109
rect 28 107 30 109
rect 24 105 30 107
rect 40 110 49 112
rect 40 108 42 110
rect 44 108 49 110
rect 40 106 49 108
rect 14 103 20 105
rect 14 100 16 103
rect 27 100 29 105
rect 47 100 49 106
rect 55 110 61 112
rect 69 111 71 115
rect 79 112 81 115
rect 90 112 92 115
rect 55 108 57 110
rect 59 108 61 110
rect 55 107 61 108
rect 77 110 83 112
rect 77 108 79 110
rect 81 108 83 110
rect 55 105 69 107
rect 67 102 69 105
rect 77 106 83 108
rect 88 110 94 112
rect 88 108 90 110
rect 92 108 94 110
rect 88 106 94 108
rect 114 109 116 123
rect 214 133 216 145
rect 245 137 247 141
rect 259 137 261 141
rect 269 137 271 145
rect 279 137 281 142
rect 314 145 371 147
rect 190 128 192 133
rect 227 128 229 133
rect 127 111 129 115
rect 145 112 147 115
rect 159 112 161 115
rect 125 109 131 111
rect 114 107 120 109
rect 77 102 79 106
rect 88 102 90 106
rect 114 105 116 107
rect 118 105 120 107
rect 125 107 127 109
rect 129 107 131 109
rect 125 105 131 107
rect 140 110 149 112
rect 140 108 142 110
rect 144 108 149 110
rect 140 106 149 108
rect 114 103 120 105
rect 14 81 16 93
rect 27 85 29 90
rect 57 97 59 101
rect 47 85 49 89
rect 114 100 116 103
rect 127 100 129 105
rect 147 100 149 106
rect 155 110 161 112
rect 169 111 171 115
rect 179 112 181 115
rect 190 112 192 115
rect 155 108 157 110
rect 159 108 161 110
rect 155 107 161 108
rect 177 110 183 112
rect 177 108 179 110
rect 181 108 183 110
rect 155 105 169 107
rect 167 102 169 105
rect 177 106 183 108
rect 188 110 194 112
rect 188 108 190 110
rect 192 108 194 110
rect 188 106 194 108
rect 214 109 216 123
rect 314 133 316 145
rect 345 137 347 141
rect 359 137 361 141
rect 369 137 371 145
rect 379 137 381 142
rect 416 145 473 147
rect 290 128 292 133
rect 327 128 329 133
rect 227 111 229 115
rect 245 112 247 115
rect 259 112 261 115
rect 224 109 230 111
rect 214 107 220 109
rect 177 102 179 106
rect 188 102 190 106
rect 214 105 216 107
rect 218 105 220 107
rect 224 107 226 109
rect 228 107 230 109
rect 224 105 230 107
rect 240 110 249 112
rect 240 108 242 110
rect 244 108 249 110
rect 240 106 249 108
rect 214 103 220 105
rect 67 86 69 91
rect 77 86 79 91
rect 88 88 90 92
rect 57 81 59 86
rect 14 79 59 81
rect 114 81 116 93
rect 127 85 129 90
rect 157 97 159 101
rect 147 85 149 89
rect 214 100 216 103
rect 227 100 229 105
rect 247 100 249 106
rect 255 110 261 112
rect 269 111 271 115
rect 279 112 281 115
rect 290 112 292 115
rect 255 108 257 110
rect 259 108 261 110
rect 255 107 261 108
rect 277 110 283 112
rect 277 108 279 110
rect 281 108 283 110
rect 255 105 269 107
rect 267 102 269 105
rect 277 106 283 108
rect 288 110 294 112
rect 288 108 290 110
rect 292 108 294 110
rect 288 106 294 108
rect 314 109 316 123
rect 416 133 418 145
rect 447 137 449 141
rect 461 137 463 141
rect 471 137 473 145
rect 481 137 483 142
rect 516 145 573 147
rect 390 128 392 133
rect 429 128 431 133
rect 327 111 329 115
rect 345 112 347 115
rect 359 112 361 115
rect 324 109 330 111
rect 314 107 320 109
rect 277 102 279 106
rect 288 102 290 106
rect 314 105 316 107
rect 318 105 320 107
rect 324 107 326 109
rect 328 107 330 109
rect 324 105 330 107
rect 340 110 349 112
rect 340 108 342 110
rect 344 108 349 110
rect 340 106 349 108
rect 314 103 320 105
rect 167 86 169 91
rect 177 86 179 91
rect 188 88 190 92
rect 157 81 159 86
rect 114 79 159 81
rect 214 81 216 93
rect 227 85 229 90
rect 257 97 259 101
rect 247 85 249 89
rect 314 100 316 103
rect 327 100 329 105
rect 347 100 349 106
rect 355 110 361 112
rect 369 111 371 115
rect 379 112 381 115
rect 390 112 392 115
rect 355 108 357 110
rect 359 108 361 110
rect 355 107 361 108
rect 377 110 383 112
rect 377 108 379 110
rect 381 108 383 110
rect 355 105 369 107
rect 367 102 369 105
rect 377 106 383 108
rect 388 110 394 112
rect 388 108 390 110
rect 392 108 394 110
rect 388 106 394 108
rect 416 109 418 123
rect 516 133 518 145
rect 547 137 549 141
rect 561 137 563 141
rect 571 137 573 145
rect 581 137 583 142
rect 616 145 673 147
rect 492 128 494 133
rect 529 128 531 133
rect 429 111 431 115
rect 447 112 449 115
rect 461 112 463 115
rect 426 109 432 111
rect 416 107 422 109
rect 377 102 379 106
rect 388 102 390 106
rect 416 105 418 107
rect 420 105 422 107
rect 426 107 428 109
rect 430 107 432 109
rect 426 105 432 107
rect 442 110 451 112
rect 442 108 444 110
rect 446 108 451 110
rect 442 106 451 108
rect 416 103 422 105
rect 267 86 269 91
rect 277 86 279 91
rect 288 88 290 92
rect 257 81 259 86
rect 214 79 259 81
rect 314 81 316 93
rect 327 85 329 90
rect 357 97 359 101
rect 347 85 349 89
rect 416 100 418 103
rect 429 100 431 105
rect 449 100 451 106
rect 457 110 463 112
rect 471 111 473 115
rect 481 112 483 115
rect 492 112 494 115
rect 457 108 459 110
rect 461 108 463 110
rect 457 107 463 108
rect 479 110 485 112
rect 479 108 481 110
rect 483 108 485 110
rect 457 105 471 107
rect 469 102 471 105
rect 479 106 485 108
rect 490 110 496 112
rect 490 108 492 110
rect 494 108 496 110
rect 490 106 496 108
rect 516 109 518 123
rect 616 133 618 145
rect 647 137 649 141
rect 661 137 663 141
rect 671 137 673 145
rect 681 137 683 142
rect 716 145 773 147
rect 592 128 594 133
rect 629 128 631 133
rect 529 111 531 115
rect 547 112 549 115
rect 561 112 563 115
rect 526 109 532 111
rect 516 107 522 109
rect 479 102 481 106
rect 490 102 492 106
rect 516 105 518 107
rect 520 105 522 107
rect 526 107 528 109
rect 530 107 532 109
rect 526 105 532 107
rect 542 110 551 112
rect 542 108 544 110
rect 546 108 551 110
rect 542 106 551 108
rect 516 103 522 105
rect 367 86 369 91
rect 377 86 379 91
rect 388 88 390 92
rect 357 81 359 86
rect 314 79 359 81
rect 416 81 418 93
rect 429 85 431 90
rect 459 97 461 101
rect 449 85 451 89
rect 516 100 518 103
rect 529 100 531 105
rect 549 100 551 106
rect 557 110 563 112
rect 571 111 573 115
rect 581 112 583 115
rect 592 112 594 115
rect 557 108 559 110
rect 561 108 563 110
rect 557 107 563 108
rect 579 110 585 112
rect 579 108 581 110
rect 583 108 585 110
rect 557 105 571 107
rect 569 102 571 105
rect 579 106 585 108
rect 590 110 596 112
rect 590 108 592 110
rect 594 108 596 110
rect 590 106 596 108
rect 616 109 618 123
rect 716 133 718 145
rect 747 137 749 141
rect 761 137 763 141
rect 771 137 773 145
rect 781 137 783 142
rect 692 128 694 133
rect 729 128 731 133
rect 629 111 631 115
rect 647 112 649 115
rect 661 112 663 115
rect 626 109 632 111
rect 616 107 622 109
rect 579 102 581 106
rect 590 102 592 106
rect 616 105 618 107
rect 620 105 622 107
rect 626 107 628 109
rect 630 107 632 109
rect 626 105 632 107
rect 642 110 651 112
rect 642 108 644 110
rect 646 108 651 110
rect 642 106 651 108
rect 616 103 622 105
rect 469 86 471 91
rect 479 86 481 91
rect 490 88 492 92
rect 459 81 461 86
rect 416 79 461 81
rect 516 81 518 93
rect 529 85 531 90
rect 559 97 561 101
rect 549 85 551 89
rect 616 100 618 103
rect 629 100 631 105
rect 649 100 651 106
rect 657 110 663 112
rect 671 111 673 115
rect 681 112 683 115
rect 692 112 694 115
rect 657 108 659 110
rect 661 108 663 110
rect 657 107 663 108
rect 679 110 685 112
rect 679 108 681 110
rect 683 108 685 110
rect 657 105 671 107
rect 669 102 671 105
rect 679 106 685 108
rect 690 110 696 112
rect 690 108 692 110
rect 694 108 696 110
rect 690 106 696 108
rect 716 109 718 123
rect 792 128 794 133
rect 729 111 731 115
rect 747 112 749 115
rect 761 112 763 115
rect 726 109 732 111
rect 716 107 722 109
rect 679 102 681 106
rect 690 102 692 106
rect 716 105 718 107
rect 720 105 722 107
rect 726 107 728 109
rect 730 107 732 109
rect 726 105 732 107
rect 742 110 751 112
rect 742 108 744 110
rect 746 108 751 110
rect 742 106 751 108
rect 716 103 722 105
rect 569 86 571 91
rect 579 86 581 91
rect 590 88 592 92
rect 559 81 561 86
rect 516 79 561 81
rect 616 81 618 93
rect 629 85 631 90
rect 659 97 661 101
rect 649 85 651 89
rect 716 100 718 103
rect 729 100 731 105
rect 749 100 751 106
rect 757 110 763 112
rect 771 111 773 115
rect 781 112 783 115
rect 792 112 794 115
rect 757 108 759 110
rect 761 108 763 110
rect 757 107 763 108
rect 779 110 785 112
rect 779 108 781 110
rect 783 108 785 110
rect 757 105 771 107
rect 769 102 771 105
rect 779 106 785 108
rect 790 110 796 112
rect 790 108 792 110
rect 794 108 796 110
rect 790 106 796 108
rect 779 102 781 106
rect 790 102 792 106
rect 669 86 671 91
rect 679 86 681 91
rect 690 88 692 92
rect 659 81 661 86
rect 616 79 661 81
rect 716 81 718 93
rect 729 85 731 90
rect 759 97 761 101
rect 749 85 751 89
rect 769 86 771 91
rect 779 86 781 91
rect 790 88 792 92
rect 759 81 761 86
rect 716 79 761 81
rect 47 73 92 75
rect 47 68 49 73
rect 16 62 18 66
rect 27 63 29 68
rect 37 63 39 68
rect 57 65 59 69
rect 47 53 49 57
rect 77 64 79 69
rect 90 61 92 73
rect 147 73 192 75
rect 147 68 149 73
rect 116 62 118 66
rect 127 63 129 68
rect 137 63 139 68
rect 16 48 18 52
rect 27 48 29 52
rect 12 46 18 48
rect 12 44 14 46
rect 16 44 18 46
rect 12 42 18 44
rect 23 46 29 48
rect 37 49 39 52
rect 37 47 51 49
rect 23 44 25 46
rect 27 44 29 46
rect 23 42 29 44
rect 45 46 51 47
rect 45 44 47 46
rect 49 44 51 46
rect 14 39 16 42
rect 25 39 27 42
rect 35 39 37 43
rect 45 42 51 44
rect 57 48 59 54
rect 77 49 79 54
rect 90 51 92 54
rect 157 65 159 69
rect 147 53 149 57
rect 177 64 179 69
rect 190 61 192 73
rect 247 73 292 75
rect 247 68 249 73
rect 216 62 218 66
rect 227 63 229 68
rect 237 63 239 68
rect 86 49 92 51
rect 57 46 66 48
rect 57 44 62 46
rect 64 44 66 46
rect 57 42 66 44
rect 76 47 82 49
rect 76 45 78 47
rect 80 45 82 47
rect 86 47 88 49
rect 90 47 92 49
rect 116 48 118 52
rect 127 48 129 52
rect 86 45 92 47
rect 76 43 82 45
rect 45 39 47 42
rect 59 39 61 42
rect 77 39 79 43
rect 14 21 16 26
rect 90 31 92 45
rect 112 46 118 48
rect 112 44 114 46
rect 116 44 118 46
rect 112 42 118 44
rect 123 46 129 48
rect 137 49 139 52
rect 137 47 151 49
rect 123 44 125 46
rect 127 44 129 46
rect 123 42 129 44
rect 145 46 151 47
rect 145 44 147 46
rect 149 44 151 46
rect 114 39 116 42
rect 125 39 127 42
rect 135 39 137 43
rect 145 42 151 44
rect 157 48 159 54
rect 177 49 179 54
rect 190 51 192 54
rect 257 65 259 69
rect 247 53 249 57
rect 277 64 279 69
rect 290 61 292 73
rect 347 73 392 75
rect 347 68 349 73
rect 316 62 318 66
rect 327 63 329 68
rect 337 63 339 68
rect 186 49 192 51
rect 157 46 166 48
rect 157 44 162 46
rect 164 44 166 46
rect 157 42 166 44
rect 176 47 182 49
rect 176 45 178 47
rect 180 45 182 47
rect 186 47 188 49
rect 190 47 192 49
rect 216 48 218 52
rect 227 48 229 52
rect 186 45 192 47
rect 176 43 182 45
rect 145 39 147 42
rect 159 39 161 42
rect 177 39 179 43
rect 77 21 79 26
rect 114 21 116 26
rect 25 12 27 17
rect 35 9 37 17
rect 45 13 47 17
rect 59 13 61 17
rect 90 9 92 21
rect 190 31 192 45
rect 212 46 218 48
rect 212 44 214 46
rect 216 44 218 46
rect 212 42 218 44
rect 223 46 229 48
rect 237 49 239 52
rect 237 47 251 49
rect 223 44 225 46
rect 227 44 229 46
rect 223 42 229 44
rect 245 46 251 47
rect 245 44 247 46
rect 249 44 251 46
rect 214 39 216 42
rect 225 39 227 42
rect 235 39 237 43
rect 245 42 251 44
rect 257 48 259 54
rect 277 49 279 54
rect 290 51 292 54
rect 357 65 359 69
rect 347 53 349 57
rect 377 64 379 69
rect 390 61 392 73
rect 447 73 492 75
rect 447 68 449 73
rect 416 62 418 66
rect 427 63 429 68
rect 437 63 439 68
rect 286 49 292 51
rect 257 46 266 48
rect 257 44 262 46
rect 264 44 266 46
rect 257 42 266 44
rect 276 47 282 49
rect 276 45 278 47
rect 280 45 282 47
rect 286 47 288 49
rect 290 47 292 49
rect 316 48 318 52
rect 327 48 329 52
rect 286 45 292 47
rect 276 43 282 45
rect 245 39 247 42
rect 259 39 261 42
rect 277 39 279 43
rect 177 21 179 26
rect 214 21 216 26
rect 35 7 92 9
rect 125 12 127 17
rect 135 9 137 17
rect 145 13 147 17
rect 159 13 161 17
rect 190 9 192 21
rect 290 31 292 45
rect 312 46 318 48
rect 312 44 314 46
rect 316 44 318 46
rect 312 42 318 44
rect 323 46 329 48
rect 337 49 339 52
rect 337 47 351 49
rect 323 44 325 46
rect 327 44 329 46
rect 323 42 329 44
rect 345 46 351 47
rect 345 44 347 46
rect 349 44 351 46
rect 314 39 316 42
rect 325 39 327 42
rect 335 39 337 43
rect 345 42 351 44
rect 357 48 359 54
rect 377 49 379 54
rect 390 51 392 54
rect 457 65 459 69
rect 447 53 449 57
rect 477 64 479 69
rect 490 61 492 73
rect 547 73 592 75
rect 547 68 549 73
rect 516 62 518 66
rect 527 63 529 68
rect 537 63 539 68
rect 386 49 392 51
rect 357 46 366 48
rect 357 44 362 46
rect 364 44 366 46
rect 357 42 366 44
rect 376 47 382 49
rect 376 45 378 47
rect 380 45 382 47
rect 386 47 388 49
rect 390 47 392 49
rect 416 48 418 52
rect 427 48 429 52
rect 386 45 392 47
rect 376 43 382 45
rect 345 39 347 42
rect 359 39 361 42
rect 377 39 379 43
rect 277 21 279 26
rect 314 21 316 26
rect 135 7 192 9
rect 225 12 227 17
rect 235 9 237 17
rect 245 13 247 17
rect 259 13 261 17
rect 290 9 292 21
rect 390 31 392 45
rect 412 46 418 48
rect 412 44 414 46
rect 416 44 418 46
rect 412 42 418 44
rect 423 46 429 48
rect 437 49 439 52
rect 437 47 451 49
rect 423 44 425 46
rect 427 44 429 46
rect 423 42 429 44
rect 445 46 451 47
rect 445 44 447 46
rect 449 44 451 46
rect 414 39 416 42
rect 425 39 427 42
rect 435 39 437 43
rect 445 42 451 44
rect 457 48 459 54
rect 477 49 479 54
rect 490 51 492 54
rect 557 65 559 69
rect 547 53 549 57
rect 577 64 579 69
rect 590 61 592 73
rect 647 73 692 75
rect 647 68 649 73
rect 616 62 618 66
rect 627 63 629 68
rect 637 63 639 68
rect 486 49 492 51
rect 457 46 466 48
rect 457 44 462 46
rect 464 44 466 46
rect 457 42 466 44
rect 476 47 482 49
rect 476 45 478 47
rect 480 45 482 47
rect 486 47 488 49
rect 490 47 492 49
rect 516 48 518 52
rect 527 48 529 52
rect 486 45 492 47
rect 476 43 482 45
rect 445 39 447 42
rect 459 39 461 42
rect 477 39 479 43
rect 377 21 379 26
rect 414 21 416 26
rect 235 7 292 9
rect 325 12 327 17
rect 335 9 337 17
rect 345 13 347 17
rect 359 13 361 17
rect 390 9 392 21
rect 490 31 492 45
rect 512 46 518 48
rect 512 44 514 46
rect 516 44 518 46
rect 512 42 518 44
rect 523 46 529 48
rect 537 49 539 52
rect 537 47 551 49
rect 523 44 525 46
rect 527 44 529 46
rect 523 42 529 44
rect 545 46 551 47
rect 545 44 547 46
rect 549 44 551 46
rect 514 39 516 42
rect 525 39 527 42
rect 535 39 537 43
rect 545 42 551 44
rect 557 48 559 54
rect 577 49 579 54
rect 590 51 592 54
rect 657 65 659 69
rect 647 53 649 57
rect 677 64 679 69
rect 690 61 692 73
rect 747 73 792 75
rect 747 68 749 73
rect 716 62 718 66
rect 727 63 729 68
rect 737 63 739 68
rect 586 49 592 51
rect 557 46 566 48
rect 557 44 562 46
rect 564 44 566 46
rect 557 42 566 44
rect 576 47 582 49
rect 576 45 578 47
rect 580 45 582 47
rect 586 47 588 49
rect 590 47 592 49
rect 616 48 618 52
rect 627 48 629 52
rect 586 45 592 47
rect 576 43 582 45
rect 545 39 547 42
rect 559 39 561 42
rect 577 39 579 43
rect 477 21 479 26
rect 514 21 516 26
rect 335 7 392 9
rect 425 12 427 17
rect 435 9 437 17
rect 445 13 447 17
rect 459 13 461 17
rect 490 9 492 21
rect 590 31 592 45
rect 612 46 618 48
rect 612 44 614 46
rect 616 44 618 46
rect 612 42 618 44
rect 623 46 629 48
rect 637 49 639 52
rect 637 47 651 49
rect 623 44 625 46
rect 627 44 629 46
rect 623 42 629 44
rect 645 46 651 47
rect 645 44 647 46
rect 649 44 651 46
rect 614 39 616 42
rect 625 39 627 42
rect 635 39 637 43
rect 645 42 651 44
rect 657 48 659 54
rect 677 49 679 54
rect 690 51 692 54
rect 757 65 759 69
rect 747 53 749 57
rect 777 64 779 69
rect 790 61 792 73
rect 686 49 692 51
rect 657 46 666 48
rect 657 44 662 46
rect 664 44 666 46
rect 657 42 666 44
rect 676 47 682 49
rect 676 45 678 47
rect 680 45 682 47
rect 686 47 688 49
rect 690 47 692 49
rect 716 48 718 52
rect 727 48 729 52
rect 686 45 692 47
rect 676 43 682 45
rect 645 39 647 42
rect 659 39 661 42
rect 677 39 679 43
rect 577 21 579 26
rect 614 21 616 26
rect 435 7 492 9
rect 525 12 527 17
rect 535 9 537 17
rect 545 13 547 17
rect 559 13 561 17
rect 590 9 592 21
rect 690 31 692 45
rect 712 46 718 48
rect 712 44 714 46
rect 716 44 718 46
rect 712 42 718 44
rect 723 46 729 48
rect 737 49 739 52
rect 737 47 751 49
rect 723 44 725 46
rect 727 44 729 46
rect 723 42 729 44
rect 745 46 751 47
rect 745 44 747 46
rect 749 44 751 46
rect 714 39 716 42
rect 725 39 727 42
rect 735 39 737 43
rect 745 42 751 44
rect 757 48 759 54
rect 777 49 779 54
rect 790 51 792 54
rect 786 49 792 51
rect 757 46 766 48
rect 757 44 762 46
rect 764 44 766 46
rect 757 42 766 44
rect 776 47 782 49
rect 776 45 778 47
rect 780 45 782 47
rect 786 47 788 49
rect 790 47 792 49
rect 786 45 792 47
rect 776 43 782 45
rect 745 39 747 42
rect 759 39 761 42
rect 777 39 779 43
rect 677 21 679 26
rect 714 21 716 26
rect 535 7 592 9
rect 625 12 627 17
rect 635 9 637 17
rect 645 13 647 17
rect 659 13 661 17
rect 690 9 692 21
rect 790 31 792 45
rect 777 21 779 26
rect 635 7 692 9
rect 725 12 727 17
rect 735 9 737 17
rect 745 13 747 17
rect 759 13 761 17
rect 790 9 792 21
rect 735 7 792 9
<< ndif >>
rect 82 357 88 359
rect 42 351 47 356
rect 20 350 27 351
rect 11 346 16 350
rect 9 344 16 346
rect 9 342 11 344
rect 13 342 16 344
rect 9 340 16 342
rect 18 349 27 350
rect 18 347 22 349
rect 24 347 27 349
rect 18 340 27 347
rect 29 344 37 351
rect 29 342 32 344
rect 34 342 37 344
rect 29 340 37 342
rect 39 349 47 351
rect 39 347 42 349
rect 44 347 47 349
rect 39 345 47 347
rect 49 353 54 356
rect 49 349 57 353
rect 49 347 52 349
rect 54 347 57 349
rect 49 345 57 347
rect 39 340 44 345
rect 52 342 57 345
rect 59 351 66 353
rect 82 355 84 357
rect 86 355 88 357
rect 82 352 88 355
rect 59 349 62 351
rect 64 349 66 351
rect 59 342 66 349
rect 72 348 77 352
rect 70 346 77 348
rect 70 344 72 346
rect 74 344 77 346
rect 70 342 77 344
rect 79 349 88 352
rect 182 357 188 359
rect 142 351 147 356
rect 120 350 127 351
rect 79 342 90 349
rect 92 346 99 349
rect 111 346 116 350
rect 92 344 95 346
rect 97 344 99 346
rect 92 342 99 344
rect 109 344 116 346
rect 109 342 111 344
rect 113 342 116 344
rect 109 340 116 342
rect 118 349 127 350
rect 118 347 122 349
rect 124 347 127 349
rect 118 340 127 347
rect 129 344 137 351
rect 129 342 132 344
rect 134 342 137 344
rect 129 340 137 342
rect 139 349 147 351
rect 139 347 142 349
rect 144 347 147 349
rect 139 345 147 347
rect 149 353 154 356
rect 149 349 157 353
rect 149 347 152 349
rect 154 347 157 349
rect 149 345 157 347
rect 139 340 144 345
rect 152 342 157 345
rect 159 351 166 353
rect 182 355 184 357
rect 186 355 188 357
rect 182 352 188 355
rect 159 349 162 351
rect 164 349 166 351
rect 159 342 166 349
rect 172 348 177 352
rect 170 346 177 348
rect 170 344 172 346
rect 174 344 177 346
rect 170 342 177 344
rect 179 349 188 352
rect 282 357 288 359
rect 242 351 247 356
rect 220 350 227 351
rect 179 342 190 349
rect 192 346 199 349
rect 211 346 216 350
rect 192 344 195 346
rect 197 344 199 346
rect 192 342 199 344
rect 209 344 216 346
rect 209 342 211 344
rect 213 342 216 344
rect 209 340 216 342
rect 218 349 227 350
rect 218 347 222 349
rect 224 347 227 349
rect 218 340 227 347
rect 229 344 237 351
rect 229 342 232 344
rect 234 342 237 344
rect 229 340 237 342
rect 239 349 247 351
rect 239 347 242 349
rect 244 347 247 349
rect 239 345 247 347
rect 249 353 254 356
rect 249 349 257 353
rect 249 347 252 349
rect 254 347 257 349
rect 249 345 257 347
rect 239 340 244 345
rect 252 342 257 345
rect 259 351 266 353
rect 282 355 284 357
rect 286 355 288 357
rect 282 352 288 355
rect 259 349 262 351
rect 264 349 266 351
rect 259 342 266 349
rect 272 348 277 352
rect 270 346 277 348
rect 270 344 272 346
rect 274 344 277 346
rect 270 342 277 344
rect 279 349 288 352
rect 382 357 388 359
rect 342 351 347 356
rect 320 350 327 351
rect 279 342 290 349
rect 292 346 299 349
rect 311 346 316 350
rect 292 344 295 346
rect 297 344 299 346
rect 292 342 299 344
rect 309 344 316 346
rect 309 342 311 344
rect 313 342 316 344
rect 309 340 316 342
rect 318 349 327 350
rect 318 347 322 349
rect 324 347 327 349
rect 318 340 327 347
rect 329 344 337 351
rect 329 342 332 344
rect 334 342 337 344
rect 329 340 337 342
rect 339 349 347 351
rect 339 347 342 349
rect 344 347 347 349
rect 339 345 347 347
rect 349 353 354 356
rect 349 349 357 353
rect 349 347 352 349
rect 354 347 357 349
rect 349 345 357 347
rect 339 340 344 345
rect 352 342 357 345
rect 359 351 366 353
rect 382 355 384 357
rect 386 355 388 357
rect 382 352 388 355
rect 359 349 362 351
rect 364 349 366 351
rect 359 342 366 349
rect 372 348 377 352
rect 370 346 377 348
rect 370 344 372 346
rect 374 344 377 346
rect 370 342 377 344
rect 379 349 388 352
rect 482 357 488 359
rect 442 351 447 356
rect 420 350 427 351
rect 379 342 390 349
rect 392 346 399 349
rect 411 346 416 350
rect 392 344 395 346
rect 397 344 399 346
rect 392 342 399 344
rect 409 344 416 346
rect 409 342 411 344
rect 413 342 416 344
rect 409 340 416 342
rect 418 349 427 350
rect 418 347 422 349
rect 424 347 427 349
rect 418 340 427 347
rect 429 344 437 351
rect 429 342 432 344
rect 434 342 437 344
rect 429 340 437 342
rect 439 349 447 351
rect 439 347 442 349
rect 444 347 447 349
rect 439 345 447 347
rect 449 353 454 356
rect 449 349 457 353
rect 449 347 452 349
rect 454 347 457 349
rect 449 345 457 347
rect 439 340 444 345
rect 452 342 457 345
rect 459 351 466 353
rect 482 355 484 357
rect 486 355 488 357
rect 482 352 488 355
rect 459 349 462 351
rect 464 349 466 351
rect 459 342 466 349
rect 472 348 477 352
rect 470 346 477 348
rect 470 344 472 346
rect 474 344 477 346
rect 470 342 477 344
rect 479 349 488 352
rect 582 357 588 359
rect 542 351 547 356
rect 520 350 527 351
rect 479 342 490 349
rect 492 346 499 349
rect 511 346 516 350
rect 492 344 495 346
rect 497 344 499 346
rect 492 342 499 344
rect 509 344 516 346
rect 509 342 511 344
rect 513 342 516 344
rect 509 340 516 342
rect 518 349 527 350
rect 518 347 522 349
rect 524 347 527 349
rect 518 340 527 347
rect 529 344 537 351
rect 529 342 532 344
rect 534 342 537 344
rect 529 340 537 342
rect 539 349 547 351
rect 539 347 542 349
rect 544 347 547 349
rect 539 345 547 347
rect 549 353 554 356
rect 549 349 557 353
rect 549 347 552 349
rect 554 347 557 349
rect 549 345 557 347
rect 539 340 544 345
rect 552 342 557 345
rect 559 351 566 353
rect 582 355 584 357
rect 586 355 588 357
rect 582 352 588 355
rect 559 349 562 351
rect 564 349 566 351
rect 559 342 566 349
rect 572 348 577 352
rect 570 346 577 348
rect 570 344 572 346
rect 574 344 577 346
rect 570 342 577 344
rect 579 349 588 352
rect 682 357 688 359
rect 642 351 647 356
rect 620 350 627 351
rect 579 342 590 349
rect 592 346 599 349
rect 611 346 616 350
rect 592 344 595 346
rect 597 344 599 346
rect 592 342 599 344
rect 609 344 616 346
rect 609 342 611 344
rect 613 342 616 344
rect 609 340 616 342
rect 618 349 627 350
rect 618 347 622 349
rect 624 347 627 349
rect 618 340 627 347
rect 629 344 637 351
rect 629 342 632 344
rect 634 342 637 344
rect 629 340 637 342
rect 639 349 647 351
rect 639 347 642 349
rect 644 347 647 349
rect 639 345 647 347
rect 649 353 654 356
rect 649 349 657 353
rect 649 347 652 349
rect 654 347 657 349
rect 649 345 657 347
rect 639 340 644 345
rect 652 342 657 345
rect 659 351 666 353
rect 682 355 684 357
rect 686 355 688 357
rect 682 352 688 355
rect 659 349 662 351
rect 664 349 666 351
rect 659 342 666 349
rect 672 348 677 352
rect 670 346 677 348
rect 670 344 672 346
rect 674 344 677 346
rect 670 342 677 344
rect 679 349 688 352
rect 782 357 788 359
rect 742 351 747 356
rect 720 350 727 351
rect 679 342 690 349
rect 692 346 699 349
rect 711 346 716 350
rect 692 344 695 346
rect 697 344 699 346
rect 692 342 699 344
rect 709 344 716 346
rect 709 342 711 344
rect 713 342 716 344
rect 709 340 716 342
rect 718 349 727 350
rect 718 347 722 349
rect 724 347 727 349
rect 718 340 727 347
rect 729 344 737 351
rect 729 342 732 344
rect 734 342 737 344
rect 729 340 737 342
rect 739 349 747 351
rect 739 347 742 349
rect 744 347 747 349
rect 739 345 747 347
rect 749 353 754 356
rect 749 349 757 353
rect 749 347 752 349
rect 754 347 757 349
rect 749 345 757 347
rect 739 340 744 345
rect 752 342 757 345
rect 759 351 766 353
rect 782 355 784 357
rect 786 355 788 357
rect 782 352 788 355
rect 759 349 762 351
rect 764 349 766 351
rect 759 342 766 349
rect 772 348 777 352
rect 770 346 777 348
rect 770 344 772 346
rect 774 344 777 346
rect 770 342 777 344
rect 779 349 788 352
rect 779 342 790 349
rect 792 346 799 349
rect 792 344 795 346
rect 797 344 799 346
rect 792 342 799 344
rect 7 242 14 244
rect 7 240 9 242
rect 11 240 14 242
rect 7 237 14 240
rect 16 237 27 244
rect 18 234 27 237
rect 29 242 36 244
rect 29 240 32 242
rect 34 240 36 242
rect 29 238 36 240
rect 29 234 34 238
rect 40 237 47 244
rect 40 235 42 237
rect 44 235 47 237
rect 18 231 24 234
rect 18 229 20 231
rect 22 229 24 231
rect 40 233 47 235
rect 49 241 54 244
rect 62 241 67 246
rect 49 239 57 241
rect 49 237 52 239
rect 54 237 57 239
rect 49 233 57 237
rect 52 230 57 233
rect 59 239 67 241
rect 59 237 62 239
rect 64 237 67 239
rect 59 235 67 237
rect 69 244 77 246
rect 69 242 72 244
rect 74 242 77 244
rect 69 235 77 242
rect 79 239 88 246
rect 79 237 82 239
rect 84 237 88 239
rect 79 236 88 237
rect 90 244 97 246
rect 90 242 93 244
rect 95 242 97 244
rect 90 240 97 242
rect 107 242 114 244
rect 107 240 109 242
rect 111 240 114 242
rect 90 236 95 240
rect 107 237 114 240
rect 116 237 127 244
rect 79 235 86 236
rect 59 230 64 235
rect 18 227 24 229
rect 118 234 127 237
rect 129 242 136 244
rect 129 240 132 242
rect 134 240 136 242
rect 129 238 136 240
rect 129 234 134 238
rect 140 237 147 244
rect 140 235 142 237
rect 144 235 147 237
rect 118 231 124 234
rect 118 229 120 231
rect 122 229 124 231
rect 140 233 147 235
rect 149 241 154 244
rect 162 241 167 246
rect 149 239 157 241
rect 149 237 152 239
rect 154 237 157 239
rect 149 233 157 237
rect 152 230 157 233
rect 159 239 167 241
rect 159 237 162 239
rect 164 237 167 239
rect 159 235 167 237
rect 169 244 177 246
rect 169 242 172 244
rect 174 242 177 244
rect 169 235 177 242
rect 179 239 188 246
rect 179 237 182 239
rect 184 237 188 239
rect 179 236 188 237
rect 190 244 197 246
rect 190 242 193 244
rect 195 242 197 244
rect 190 240 197 242
rect 207 242 214 244
rect 207 240 209 242
rect 211 240 214 242
rect 190 236 195 240
rect 207 237 214 240
rect 216 237 227 244
rect 179 235 186 236
rect 159 230 164 235
rect 118 227 124 229
rect 218 234 227 237
rect 229 242 236 244
rect 229 240 232 242
rect 234 240 236 242
rect 229 238 236 240
rect 229 234 234 238
rect 240 237 247 244
rect 240 235 242 237
rect 244 235 247 237
rect 218 231 224 234
rect 218 229 220 231
rect 222 229 224 231
rect 240 233 247 235
rect 249 241 254 244
rect 262 241 267 246
rect 249 239 257 241
rect 249 237 252 239
rect 254 237 257 239
rect 249 233 257 237
rect 252 230 257 233
rect 259 239 267 241
rect 259 237 262 239
rect 264 237 267 239
rect 259 235 267 237
rect 269 244 277 246
rect 269 242 272 244
rect 274 242 277 244
rect 269 235 277 242
rect 279 239 288 246
rect 279 237 282 239
rect 284 237 288 239
rect 279 236 288 237
rect 290 244 297 246
rect 290 242 293 244
rect 295 242 297 244
rect 290 240 297 242
rect 307 242 314 244
rect 307 240 309 242
rect 311 240 314 242
rect 290 236 295 240
rect 307 237 314 240
rect 316 237 327 244
rect 279 235 286 236
rect 259 230 264 235
rect 218 227 224 229
rect 318 234 327 237
rect 329 242 336 244
rect 329 240 332 242
rect 334 240 336 242
rect 329 238 336 240
rect 329 234 334 238
rect 340 237 347 244
rect 340 235 342 237
rect 344 235 347 237
rect 318 231 324 234
rect 318 229 320 231
rect 322 229 324 231
rect 340 233 347 235
rect 349 241 354 244
rect 362 241 367 246
rect 349 239 357 241
rect 349 237 352 239
rect 354 237 357 239
rect 349 233 357 237
rect 352 230 357 233
rect 359 239 367 241
rect 359 237 362 239
rect 364 237 367 239
rect 359 235 367 237
rect 369 244 377 246
rect 369 242 372 244
rect 374 242 377 244
rect 369 235 377 242
rect 379 239 388 246
rect 379 237 382 239
rect 384 237 388 239
rect 379 236 388 237
rect 390 244 397 246
rect 390 242 393 244
rect 395 242 397 244
rect 390 240 397 242
rect 409 242 416 244
rect 409 240 411 242
rect 413 240 416 242
rect 390 236 395 240
rect 409 237 416 240
rect 418 237 429 244
rect 379 235 386 236
rect 359 230 364 235
rect 318 227 324 229
rect 420 234 429 237
rect 431 242 438 244
rect 431 240 434 242
rect 436 240 438 242
rect 431 238 438 240
rect 431 234 436 238
rect 442 237 449 244
rect 442 235 444 237
rect 446 235 449 237
rect 420 231 426 234
rect 420 229 422 231
rect 424 229 426 231
rect 442 233 449 235
rect 451 241 456 244
rect 464 241 469 246
rect 451 239 459 241
rect 451 237 454 239
rect 456 237 459 239
rect 451 233 459 237
rect 454 230 459 233
rect 461 239 469 241
rect 461 237 464 239
rect 466 237 469 239
rect 461 235 469 237
rect 471 244 479 246
rect 471 242 474 244
rect 476 242 479 244
rect 471 235 479 242
rect 481 239 490 246
rect 481 237 484 239
rect 486 237 490 239
rect 481 236 490 237
rect 492 244 499 246
rect 492 242 495 244
rect 497 242 499 244
rect 492 240 499 242
rect 509 242 516 244
rect 509 240 511 242
rect 513 240 516 242
rect 492 236 497 240
rect 509 237 516 240
rect 518 237 529 244
rect 481 235 488 236
rect 461 230 466 235
rect 420 227 426 229
rect 520 234 529 237
rect 531 242 538 244
rect 531 240 534 242
rect 536 240 538 242
rect 531 238 538 240
rect 531 234 536 238
rect 542 237 549 244
rect 542 235 544 237
rect 546 235 549 237
rect 520 231 526 234
rect 520 229 522 231
rect 524 229 526 231
rect 542 233 549 235
rect 551 241 556 244
rect 564 241 569 246
rect 551 239 559 241
rect 551 237 554 239
rect 556 237 559 239
rect 551 233 559 237
rect 554 230 559 233
rect 561 239 569 241
rect 561 237 564 239
rect 566 237 569 239
rect 561 235 569 237
rect 571 244 579 246
rect 571 242 574 244
rect 576 242 579 244
rect 571 235 579 242
rect 581 239 590 246
rect 581 237 584 239
rect 586 237 590 239
rect 581 236 590 237
rect 592 244 599 246
rect 592 242 595 244
rect 597 242 599 244
rect 592 240 599 242
rect 609 242 616 244
rect 609 240 611 242
rect 613 240 616 242
rect 592 236 597 240
rect 609 237 616 240
rect 618 237 629 244
rect 581 235 588 236
rect 561 230 566 235
rect 520 227 526 229
rect 620 234 629 237
rect 631 242 638 244
rect 631 240 634 242
rect 636 240 638 242
rect 631 238 638 240
rect 631 234 636 238
rect 642 237 649 244
rect 642 235 644 237
rect 646 235 649 237
rect 620 231 626 234
rect 620 229 622 231
rect 624 229 626 231
rect 642 233 649 235
rect 651 241 656 244
rect 664 241 669 246
rect 651 239 659 241
rect 651 237 654 239
rect 656 237 659 239
rect 651 233 659 237
rect 654 230 659 233
rect 661 239 669 241
rect 661 237 664 239
rect 666 237 669 239
rect 661 235 669 237
rect 671 244 679 246
rect 671 242 674 244
rect 676 242 679 244
rect 671 235 679 242
rect 681 239 690 246
rect 681 237 684 239
rect 686 237 690 239
rect 681 236 690 237
rect 692 244 699 246
rect 692 242 695 244
rect 697 242 699 244
rect 692 240 699 242
rect 709 242 716 244
rect 709 240 711 242
rect 713 240 716 242
rect 692 236 697 240
rect 709 237 716 240
rect 718 237 729 244
rect 681 235 688 236
rect 661 230 666 235
rect 620 227 626 229
rect 720 234 729 237
rect 731 242 738 244
rect 731 240 734 242
rect 736 240 738 242
rect 731 238 738 240
rect 731 234 736 238
rect 742 237 749 244
rect 742 235 744 237
rect 746 235 749 237
rect 720 231 726 234
rect 720 229 722 231
rect 724 229 726 231
rect 742 233 749 235
rect 751 241 756 244
rect 764 241 769 246
rect 751 239 759 241
rect 751 237 754 239
rect 756 237 759 239
rect 751 233 759 237
rect 754 230 759 233
rect 761 239 769 241
rect 761 237 764 239
rect 766 237 769 239
rect 761 235 769 237
rect 771 244 779 246
rect 771 242 774 244
rect 776 242 779 244
rect 771 235 779 242
rect 781 239 790 246
rect 781 237 784 239
rect 786 237 790 239
rect 781 236 790 237
rect 792 244 799 246
rect 792 242 795 244
rect 797 242 799 244
rect 792 240 799 242
rect 792 236 797 240
rect 781 235 788 236
rect 761 230 766 235
rect 720 227 726 229
rect 18 213 24 215
rect 18 211 20 213
rect 22 211 24 213
rect 18 208 24 211
rect 52 209 57 212
rect 18 205 27 208
rect 7 202 14 205
rect 7 200 9 202
rect 11 200 14 202
rect 7 198 14 200
rect 16 198 27 205
rect 29 204 34 208
rect 40 207 47 209
rect 40 205 42 207
rect 44 205 47 207
rect 29 202 36 204
rect 29 200 32 202
rect 34 200 36 202
rect 29 198 36 200
rect 40 198 47 205
rect 49 205 57 209
rect 49 203 52 205
rect 54 203 57 205
rect 49 201 57 203
rect 59 207 64 212
rect 59 205 67 207
rect 59 203 62 205
rect 64 203 67 205
rect 59 201 67 203
rect 49 198 54 201
rect 62 196 67 201
rect 69 200 77 207
rect 69 198 72 200
rect 74 198 77 200
rect 69 196 77 198
rect 79 206 86 207
rect 79 205 88 206
rect 79 203 82 205
rect 84 203 88 205
rect 79 196 88 203
rect 90 202 95 206
rect 118 213 124 215
rect 118 211 120 213
rect 122 211 124 213
rect 118 208 124 211
rect 152 209 157 212
rect 118 205 127 208
rect 107 202 114 205
rect 90 200 97 202
rect 90 198 93 200
rect 95 198 97 200
rect 107 200 109 202
rect 111 200 114 202
rect 107 198 114 200
rect 116 198 127 205
rect 129 204 134 208
rect 140 207 147 209
rect 140 205 142 207
rect 144 205 147 207
rect 129 202 136 204
rect 129 200 132 202
rect 134 200 136 202
rect 129 198 136 200
rect 140 198 147 205
rect 149 205 157 209
rect 149 203 152 205
rect 154 203 157 205
rect 149 201 157 203
rect 159 207 164 212
rect 159 205 167 207
rect 159 203 162 205
rect 164 203 167 205
rect 159 201 167 203
rect 149 198 154 201
rect 90 196 97 198
rect 162 196 167 201
rect 169 200 177 207
rect 169 198 172 200
rect 174 198 177 200
rect 169 196 177 198
rect 179 206 186 207
rect 179 205 188 206
rect 179 203 182 205
rect 184 203 188 205
rect 179 196 188 203
rect 190 202 195 206
rect 218 213 224 215
rect 218 211 220 213
rect 222 211 224 213
rect 218 208 224 211
rect 252 209 257 212
rect 218 205 227 208
rect 207 202 214 205
rect 190 200 197 202
rect 190 198 193 200
rect 195 198 197 200
rect 207 200 209 202
rect 211 200 214 202
rect 207 198 214 200
rect 216 198 227 205
rect 229 204 234 208
rect 240 207 247 209
rect 240 205 242 207
rect 244 205 247 207
rect 229 202 236 204
rect 229 200 232 202
rect 234 200 236 202
rect 229 198 236 200
rect 240 198 247 205
rect 249 205 257 209
rect 249 203 252 205
rect 254 203 257 205
rect 249 201 257 203
rect 259 207 264 212
rect 259 205 267 207
rect 259 203 262 205
rect 264 203 267 205
rect 259 201 267 203
rect 249 198 254 201
rect 190 196 197 198
rect 262 196 267 201
rect 269 200 277 207
rect 269 198 272 200
rect 274 198 277 200
rect 269 196 277 198
rect 279 206 286 207
rect 279 205 288 206
rect 279 203 282 205
rect 284 203 288 205
rect 279 196 288 203
rect 290 202 295 206
rect 318 213 324 215
rect 318 211 320 213
rect 322 211 324 213
rect 318 208 324 211
rect 352 209 357 212
rect 318 205 327 208
rect 307 202 314 205
rect 290 200 297 202
rect 290 198 293 200
rect 295 198 297 200
rect 307 200 309 202
rect 311 200 314 202
rect 307 198 314 200
rect 316 198 327 205
rect 329 204 334 208
rect 340 207 347 209
rect 340 205 342 207
rect 344 205 347 207
rect 329 202 336 204
rect 329 200 332 202
rect 334 200 336 202
rect 329 198 336 200
rect 340 198 347 205
rect 349 205 357 209
rect 349 203 352 205
rect 354 203 357 205
rect 349 201 357 203
rect 359 207 364 212
rect 359 205 367 207
rect 359 203 362 205
rect 364 203 367 205
rect 359 201 367 203
rect 349 198 354 201
rect 290 196 297 198
rect 362 196 367 201
rect 369 200 377 207
rect 369 198 372 200
rect 374 198 377 200
rect 369 196 377 198
rect 379 206 386 207
rect 379 205 388 206
rect 379 203 382 205
rect 384 203 388 205
rect 379 196 388 203
rect 390 202 395 206
rect 420 213 426 215
rect 420 211 422 213
rect 424 211 426 213
rect 420 208 426 211
rect 454 209 459 212
rect 420 205 429 208
rect 409 202 416 205
rect 390 200 397 202
rect 390 198 393 200
rect 395 198 397 200
rect 409 200 411 202
rect 413 200 416 202
rect 409 198 416 200
rect 418 198 429 205
rect 431 204 436 208
rect 442 207 449 209
rect 442 205 444 207
rect 446 205 449 207
rect 431 202 438 204
rect 431 200 434 202
rect 436 200 438 202
rect 431 198 438 200
rect 442 198 449 205
rect 451 205 459 209
rect 451 203 454 205
rect 456 203 459 205
rect 451 201 459 203
rect 461 207 466 212
rect 461 205 469 207
rect 461 203 464 205
rect 466 203 469 205
rect 461 201 469 203
rect 451 198 456 201
rect 390 196 397 198
rect 464 196 469 201
rect 471 200 479 207
rect 471 198 474 200
rect 476 198 479 200
rect 471 196 479 198
rect 481 206 488 207
rect 481 205 490 206
rect 481 203 484 205
rect 486 203 490 205
rect 481 196 490 203
rect 492 202 497 206
rect 520 213 526 215
rect 520 211 522 213
rect 524 211 526 213
rect 520 208 526 211
rect 554 209 559 212
rect 520 205 529 208
rect 509 202 516 205
rect 492 200 499 202
rect 492 198 495 200
rect 497 198 499 200
rect 509 200 511 202
rect 513 200 516 202
rect 509 198 516 200
rect 518 198 529 205
rect 531 204 536 208
rect 542 207 549 209
rect 542 205 544 207
rect 546 205 549 207
rect 531 202 538 204
rect 531 200 534 202
rect 536 200 538 202
rect 531 198 538 200
rect 542 198 549 205
rect 551 205 559 209
rect 551 203 554 205
rect 556 203 559 205
rect 551 201 559 203
rect 561 207 566 212
rect 561 205 569 207
rect 561 203 564 205
rect 566 203 569 205
rect 561 201 569 203
rect 551 198 556 201
rect 492 196 499 198
rect 564 196 569 201
rect 571 200 579 207
rect 571 198 574 200
rect 576 198 579 200
rect 571 196 579 198
rect 581 206 588 207
rect 581 205 590 206
rect 581 203 584 205
rect 586 203 590 205
rect 581 196 590 203
rect 592 202 597 206
rect 620 213 626 215
rect 620 211 622 213
rect 624 211 626 213
rect 620 208 626 211
rect 654 209 659 212
rect 620 205 629 208
rect 609 202 616 205
rect 592 200 599 202
rect 592 198 595 200
rect 597 198 599 200
rect 609 200 611 202
rect 613 200 616 202
rect 609 198 616 200
rect 618 198 629 205
rect 631 204 636 208
rect 642 207 649 209
rect 642 205 644 207
rect 646 205 649 207
rect 631 202 638 204
rect 631 200 634 202
rect 636 200 638 202
rect 631 198 638 200
rect 642 198 649 205
rect 651 205 659 209
rect 651 203 654 205
rect 656 203 659 205
rect 651 201 659 203
rect 661 207 666 212
rect 661 205 669 207
rect 661 203 664 205
rect 666 203 669 205
rect 661 201 669 203
rect 651 198 656 201
rect 592 196 599 198
rect 664 196 669 201
rect 671 200 679 207
rect 671 198 674 200
rect 676 198 679 200
rect 671 196 679 198
rect 681 206 688 207
rect 681 205 690 206
rect 681 203 684 205
rect 686 203 690 205
rect 681 196 690 203
rect 692 202 697 206
rect 720 213 726 215
rect 720 211 722 213
rect 724 211 726 213
rect 720 208 726 211
rect 754 209 759 212
rect 720 205 729 208
rect 709 202 716 205
rect 692 200 699 202
rect 692 198 695 200
rect 697 198 699 200
rect 709 200 711 202
rect 713 200 716 202
rect 709 198 716 200
rect 718 198 729 205
rect 731 204 736 208
rect 742 207 749 209
rect 742 205 744 207
rect 746 205 749 207
rect 731 202 738 204
rect 731 200 734 202
rect 736 200 738 202
rect 731 198 738 200
rect 742 198 749 205
rect 751 205 759 209
rect 751 203 754 205
rect 756 203 759 205
rect 751 201 759 203
rect 761 207 766 212
rect 761 205 769 207
rect 761 203 764 205
rect 766 203 769 205
rect 761 201 769 203
rect 751 198 756 201
rect 692 196 699 198
rect 764 196 769 201
rect 771 200 779 207
rect 771 198 774 200
rect 776 198 779 200
rect 771 196 779 198
rect 781 206 788 207
rect 781 205 790 206
rect 781 203 784 205
rect 786 203 790 205
rect 781 196 790 203
rect 792 202 797 206
rect 792 200 799 202
rect 792 198 795 200
rect 797 198 799 200
rect 792 196 799 198
rect 7 98 14 100
rect 7 96 9 98
rect 11 96 14 98
rect 7 93 14 96
rect 16 93 27 100
rect 18 90 27 93
rect 29 98 36 100
rect 29 96 32 98
rect 34 96 36 98
rect 29 94 36 96
rect 29 90 34 94
rect 40 93 47 100
rect 40 91 42 93
rect 44 91 47 93
rect 18 87 24 90
rect 18 85 20 87
rect 22 85 24 87
rect 40 89 47 91
rect 49 97 54 100
rect 62 97 67 102
rect 49 95 57 97
rect 49 93 52 95
rect 54 93 57 95
rect 49 89 57 93
rect 52 86 57 89
rect 59 95 67 97
rect 59 93 62 95
rect 64 93 67 95
rect 59 91 67 93
rect 69 100 77 102
rect 69 98 72 100
rect 74 98 77 100
rect 69 91 77 98
rect 79 95 88 102
rect 79 93 82 95
rect 84 93 88 95
rect 79 92 88 93
rect 90 100 97 102
rect 90 98 93 100
rect 95 98 97 100
rect 90 96 97 98
rect 107 98 114 100
rect 107 96 109 98
rect 111 96 114 98
rect 90 92 95 96
rect 107 93 114 96
rect 116 93 127 100
rect 79 91 86 92
rect 59 86 64 91
rect 18 83 24 85
rect 118 90 127 93
rect 129 98 136 100
rect 129 96 132 98
rect 134 96 136 98
rect 129 94 136 96
rect 129 90 134 94
rect 140 93 147 100
rect 140 91 142 93
rect 144 91 147 93
rect 118 87 124 90
rect 118 85 120 87
rect 122 85 124 87
rect 140 89 147 91
rect 149 97 154 100
rect 162 97 167 102
rect 149 95 157 97
rect 149 93 152 95
rect 154 93 157 95
rect 149 89 157 93
rect 152 86 157 89
rect 159 95 167 97
rect 159 93 162 95
rect 164 93 167 95
rect 159 91 167 93
rect 169 100 177 102
rect 169 98 172 100
rect 174 98 177 100
rect 169 91 177 98
rect 179 95 188 102
rect 179 93 182 95
rect 184 93 188 95
rect 179 92 188 93
rect 190 100 197 102
rect 190 98 193 100
rect 195 98 197 100
rect 190 96 197 98
rect 207 98 214 100
rect 207 96 209 98
rect 211 96 214 98
rect 190 92 195 96
rect 207 93 214 96
rect 216 93 227 100
rect 179 91 186 92
rect 159 86 164 91
rect 118 83 124 85
rect 218 90 227 93
rect 229 98 236 100
rect 229 96 232 98
rect 234 96 236 98
rect 229 94 236 96
rect 229 90 234 94
rect 240 93 247 100
rect 240 91 242 93
rect 244 91 247 93
rect 218 87 224 90
rect 218 85 220 87
rect 222 85 224 87
rect 240 89 247 91
rect 249 97 254 100
rect 262 97 267 102
rect 249 95 257 97
rect 249 93 252 95
rect 254 93 257 95
rect 249 89 257 93
rect 252 86 257 89
rect 259 95 267 97
rect 259 93 262 95
rect 264 93 267 95
rect 259 91 267 93
rect 269 100 277 102
rect 269 98 272 100
rect 274 98 277 100
rect 269 91 277 98
rect 279 95 288 102
rect 279 93 282 95
rect 284 93 288 95
rect 279 92 288 93
rect 290 100 297 102
rect 290 98 293 100
rect 295 98 297 100
rect 290 96 297 98
rect 307 98 314 100
rect 307 96 309 98
rect 311 96 314 98
rect 290 92 295 96
rect 307 93 314 96
rect 316 93 327 100
rect 279 91 286 92
rect 259 86 264 91
rect 218 83 224 85
rect 318 90 327 93
rect 329 98 336 100
rect 329 96 332 98
rect 334 96 336 98
rect 329 94 336 96
rect 329 90 334 94
rect 340 93 347 100
rect 340 91 342 93
rect 344 91 347 93
rect 318 87 324 90
rect 318 85 320 87
rect 322 85 324 87
rect 340 89 347 91
rect 349 97 354 100
rect 362 97 367 102
rect 349 95 357 97
rect 349 93 352 95
rect 354 93 357 95
rect 349 89 357 93
rect 352 86 357 89
rect 359 95 367 97
rect 359 93 362 95
rect 364 93 367 95
rect 359 91 367 93
rect 369 100 377 102
rect 369 98 372 100
rect 374 98 377 100
rect 369 91 377 98
rect 379 95 388 102
rect 379 93 382 95
rect 384 93 388 95
rect 379 92 388 93
rect 390 100 397 102
rect 390 98 393 100
rect 395 98 397 100
rect 390 96 397 98
rect 409 98 416 100
rect 409 96 411 98
rect 413 96 416 98
rect 390 92 395 96
rect 409 93 416 96
rect 418 93 429 100
rect 379 91 386 92
rect 359 86 364 91
rect 318 83 324 85
rect 420 90 429 93
rect 431 98 438 100
rect 431 96 434 98
rect 436 96 438 98
rect 431 94 438 96
rect 431 90 436 94
rect 442 93 449 100
rect 442 91 444 93
rect 446 91 449 93
rect 420 87 426 90
rect 420 85 422 87
rect 424 85 426 87
rect 442 89 449 91
rect 451 97 456 100
rect 464 97 469 102
rect 451 95 459 97
rect 451 93 454 95
rect 456 93 459 95
rect 451 89 459 93
rect 454 86 459 89
rect 461 95 469 97
rect 461 93 464 95
rect 466 93 469 95
rect 461 91 469 93
rect 471 100 479 102
rect 471 98 474 100
rect 476 98 479 100
rect 471 91 479 98
rect 481 95 490 102
rect 481 93 484 95
rect 486 93 490 95
rect 481 92 490 93
rect 492 100 499 102
rect 492 98 495 100
rect 497 98 499 100
rect 492 96 499 98
rect 509 98 516 100
rect 509 96 511 98
rect 513 96 516 98
rect 492 92 497 96
rect 509 93 516 96
rect 518 93 529 100
rect 481 91 488 92
rect 461 86 466 91
rect 420 83 426 85
rect 520 90 529 93
rect 531 98 538 100
rect 531 96 534 98
rect 536 96 538 98
rect 531 94 538 96
rect 531 90 536 94
rect 542 93 549 100
rect 542 91 544 93
rect 546 91 549 93
rect 520 87 526 90
rect 520 85 522 87
rect 524 85 526 87
rect 542 89 549 91
rect 551 97 556 100
rect 564 97 569 102
rect 551 95 559 97
rect 551 93 554 95
rect 556 93 559 95
rect 551 89 559 93
rect 554 86 559 89
rect 561 95 569 97
rect 561 93 564 95
rect 566 93 569 95
rect 561 91 569 93
rect 571 100 579 102
rect 571 98 574 100
rect 576 98 579 100
rect 571 91 579 98
rect 581 95 590 102
rect 581 93 584 95
rect 586 93 590 95
rect 581 92 590 93
rect 592 100 599 102
rect 592 98 595 100
rect 597 98 599 100
rect 592 96 599 98
rect 609 98 616 100
rect 609 96 611 98
rect 613 96 616 98
rect 592 92 597 96
rect 609 93 616 96
rect 618 93 629 100
rect 581 91 588 92
rect 561 86 566 91
rect 520 83 526 85
rect 620 90 629 93
rect 631 98 638 100
rect 631 96 634 98
rect 636 96 638 98
rect 631 94 638 96
rect 631 90 636 94
rect 642 93 649 100
rect 642 91 644 93
rect 646 91 649 93
rect 620 87 626 90
rect 620 85 622 87
rect 624 85 626 87
rect 642 89 649 91
rect 651 97 656 100
rect 664 97 669 102
rect 651 95 659 97
rect 651 93 654 95
rect 656 93 659 95
rect 651 89 659 93
rect 654 86 659 89
rect 661 95 669 97
rect 661 93 664 95
rect 666 93 669 95
rect 661 91 669 93
rect 671 100 679 102
rect 671 98 674 100
rect 676 98 679 100
rect 671 91 679 98
rect 681 95 690 102
rect 681 93 684 95
rect 686 93 690 95
rect 681 92 690 93
rect 692 100 699 102
rect 692 98 695 100
rect 697 98 699 100
rect 692 96 699 98
rect 709 98 716 100
rect 709 96 711 98
rect 713 96 716 98
rect 692 92 697 96
rect 709 93 716 96
rect 718 93 729 100
rect 681 91 688 92
rect 661 86 666 91
rect 620 83 626 85
rect 720 90 729 93
rect 731 98 738 100
rect 731 96 734 98
rect 736 96 738 98
rect 731 94 738 96
rect 731 90 736 94
rect 742 93 749 100
rect 742 91 744 93
rect 746 91 749 93
rect 720 87 726 90
rect 720 85 722 87
rect 724 85 726 87
rect 742 89 749 91
rect 751 97 756 100
rect 764 97 769 102
rect 751 95 759 97
rect 751 93 754 95
rect 756 93 759 95
rect 751 89 759 93
rect 754 86 759 89
rect 761 95 769 97
rect 761 93 764 95
rect 766 93 769 95
rect 761 91 769 93
rect 771 100 779 102
rect 771 98 774 100
rect 776 98 779 100
rect 771 91 779 98
rect 781 95 790 102
rect 781 93 784 95
rect 786 93 790 95
rect 781 92 790 93
rect 792 100 799 102
rect 792 98 795 100
rect 797 98 799 100
rect 792 96 799 98
rect 792 92 797 96
rect 781 91 788 92
rect 761 86 766 91
rect 720 83 726 85
rect 82 69 88 71
rect 42 63 47 68
rect 20 62 27 63
rect 11 58 16 62
rect 9 56 16 58
rect 9 54 11 56
rect 13 54 16 56
rect 9 52 16 54
rect 18 61 27 62
rect 18 59 22 61
rect 24 59 27 61
rect 18 52 27 59
rect 29 56 37 63
rect 29 54 32 56
rect 34 54 37 56
rect 29 52 37 54
rect 39 61 47 63
rect 39 59 42 61
rect 44 59 47 61
rect 39 57 47 59
rect 49 65 54 68
rect 49 61 57 65
rect 49 59 52 61
rect 54 59 57 61
rect 49 57 57 59
rect 39 52 44 57
rect 52 54 57 57
rect 59 63 66 65
rect 82 67 84 69
rect 86 67 88 69
rect 82 64 88 67
rect 59 61 62 63
rect 64 61 66 63
rect 59 54 66 61
rect 72 60 77 64
rect 70 58 77 60
rect 70 56 72 58
rect 74 56 77 58
rect 70 54 77 56
rect 79 61 88 64
rect 182 69 188 71
rect 142 63 147 68
rect 120 62 127 63
rect 79 54 90 61
rect 92 58 99 61
rect 111 58 116 62
rect 92 56 95 58
rect 97 56 99 58
rect 92 54 99 56
rect 109 56 116 58
rect 109 54 111 56
rect 113 54 116 56
rect 109 52 116 54
rect 118 61 127 62
rect 118 59 122 61
rect 124 59 127 61
rect 118 52 127 59
rect 129 56 137 63
rect 129 54 132 56
rect 134 54 137 56
rect 129 52 137 54
rect 139 61 147 63
rect 139 59 142 61
rect 144 59 147 61
rect 139 57 147 59
rect 149 65 154 68
rect 149 61 157 65
rect 149 59 152 61
rect 154 59 157 61
rect 149 57 157 59
rect 139 52 144 57
rect 152 54 157 57
rect 159 63 166 65
rect 182 67 184 69
rect 186 67 188 69
rect 182 64 188 67
rect 159 61 162 63
rect 164 61 166 63
rect 159 54 166 61
rect 172 60 177 64
rect 170 58 177 60
rect 170 56 172 58
rect 174 56 177 58
rect 170 54 177 56
rect 179 61 188 64
rect 282 69 288 71
rect 242 63 247 68
rect 220 62 227 63
rect 179 54 190 61
rect 192 58 199 61
rect 211 58 216 62
rect 192 56 195 58
rect 197 56 199 58
rect 192 54 199 56
rect 209 56 216 58
rect 209 54 211 56
rect 213 54 216 56
rect 209 52 216 54
rect 218 61 227 62
rect 218 59 222 61
rect 224 59 227 61
rect 218 52 227 59
rect 229 56 237 63
rect 229 54 232 56
rect 234 54 237 56
rect 229 52 237 54
rect 239 61 247 63
rect 239 59 242 61
rect 244 59 247 61
rect 239 57 247 59
rect 249 65 254 68
rect 249 61 257 65
rect 249 59 252 61
rect 254 59 257 61
rect 249 57 257 59
rect 239 52 244 57
rect 252 54 257 57
rect 259 63 266 65
rect 282 67 284 69
rect 286 67 288 69
rect 282 64 288 67
rect 259 61 262 63
rect 264 61 266 63
rect 259 54 266 61
rect 272 60 277 64
rect 270 58 277 60
rect 270 56 272 58
rect 274 56 277 58
rect 270 54 277 56
rect 279 61 288 64
rect 382 69 388 71
rect 342 63 347 68
rect 320 62 327 63
rect 279 54 290 61
rect 292 58 299 61
rect 311 58 316 62
rect 292 56 295 58
rect 297 56 299 58
rect 292 54 299 56
rect 309 56 316 58
rect 309 54 311 56
rect 313 54 316 56
rect 309 52 316 54
rect 318 61 327 62
rect 318 59 322 61
rect 324 59 327 61
rect 318 52 327 59
rect 329 56 337 63
rect 329 54 332 56
rect 334 54 337 56
rect 329 52 337 54
rect 339 61 347 63
rect 339 59 342 61
rect 344 59 347 61
rect 339 57 347 59
rect 349 65 354 68
rect 349 61 357 65
rect 349 59 352 61
rect 354 59 357 61
rect 349 57 357 59
rect 339 52 344 57
rect 352 54 357 57
rect 359 63 366 65
rect 382 67 384 69
rect 386 67 388 69
rect 382 64 388 67
rect 359 61 362 63
rect 364 61 366 63
rect 359 54 366 61
rect 372 60 377 64
rect 370 58 377 60
rect 370 56 372 58
rect 374 56 377 58
rect 370 54 377 56
rect 379 61 388 64
rect 482 69 488 71
rect 442 63 447 68
rect 420 62 427 63
rect 379 54 390 61
rect 392 58 399 61
rect 411 58 416 62
rect 392 56 395 58
rect 397 56 399 58
rect 392 54 399 56
rect 409 56 416 58
rect 409 54 411 56
rect 413 54 416 56
rect 409 52 416 54
rect 418 61 427 62
rect 418 59 422 61
rect 424 59 427 61
rect 418 52 427 59
rect 429 56 437 63
rect 429 54 432 56
rect 434 54 437 56
rect 429 52 437 54
rect 439 61 447 63
rect 439 59 442 61
rect 444 59 447 61
rect 439 57 447 59
rect 449 65 454 68
rect 449 61 457 65
rect 449 59 452 61
rect 454 59 457 61
rect 449 57 457 59
rect 439 52 444 57
rect 452 54 457 57
rect 459 63 466 65
rect 482 67 484 69
rect 486 67 488 69
rect 482 64 488 67
rect 459 61 462 63
rect 464 61 466 63
rect 459 54 466 61
rect 472 60 477 64
rect 470 58 477 60
rect 470 56 472 58
rect 474 56 477 58
rect 470 54 477 56
rect 479 61 488 64
rect 582 69 588 71
rect 542 63 547 68
rect 520 62 527 63
rect 479 54 490 61
rect 492 58 499 61
rect 511 58 516 62
rect 492 56 495 58
rect 497 56 499 58
rect 492 54 499 56
rect 509 56 516 58
rect 509 54 511 56
rect 513 54 516 56
rect 509 52 516 54
rect 518 61 527 62
rect 518 59 522 61
rect 524 59 527 61
rect 518 52 527 59
rect 529 56 537 63
rect 529 54 532 56
rect 534 54 537 56
rect 529 52 537 54
rect 539 61 547 63
rect 539 59 542 61
rect 544 59 547 61
rect 539 57 547 59
rect 549 65 554 68
rect 549 61 557 65
rect 549 59 552 61
rect 554 59 557 61
rect 549 57 557 59
rect 539 52 544 57
rect 552 54 557 57
rect 559 63 566 65
rect 582 67 584 69
rect 586 67 588 69
rect 582 64 588 67
rect 559 61 562 63
rect 564 61 566 63
rect 559 54 566 61
rect 572 60 577 64
rect 570 58 577 60
rect 570 56 572 58
rect 574 56 577 58
rect 570 54 577 56
rect 579 61 588 64
rect 682 69 688 71
rect 642 63 647 68
rect 620 62 627 63
rect 579 54 590 61
rect 592 58 599 61
rect 611 58 616 62
rect 592 56 595 58
rect 597 56 599 58
rect 592 54 599 56
rect 609 56 616 58
rect 609 54 611 56
rect 613 54 616 56
rect 609 52 616 54
rect 618 61 627 62
rect 618 59 622 61
rect 624 59 627 61
rect 618 52 627 59
rect 629 56 637 63
rect 629 54 632 56
rect 634 54 637 56
rect 629 52 637 54
rect 639 61 647 63
rect 639 59 642 61
rect 644 59 647 61
rect 639 57 647 59
rect 649 65 654 68
rect 649 61 657 65
rect 649 59 652 61
rect 654 59 657 61
rect 649 57 657 59
rect 639 52 644 57
rect 652 54 657 57
rect 659 63 666 65
rect 682 67 684 69
rect 686 67 688 69
rect 682 64 688 67
rect 659 61 662 63
rect 664 61 666 63
rect 659 54 666 61
rect 672 60 677 64
rect 670 58 677 60
rect 670 56 672 58
rect 674 56 677 58
rect 670 54 677 56
rect 679 61 688 64
rect 782 69 788 71
rect 742 63 747 68
rect 720 62 727 63
rect 679 54 690 61
rect 692 58 699 61
rect 711 58 716 62
rect 692 56 695 58
rect 697 56 699 58
rect 692 54 699 56
rect 709 56 716 58
rect 709 54 711 56
rect 713 54 716 56
rect 709 52 716 54
rect 718 61 727 62
rect 718 59 722 61
rect 724 59 727 61
rect 718 52 727 59
rect 729 56 737 63
rect 729 54 732 56
rect 734 54 737 56
rect 729 52 737 54
rect 739 61 747 63
rect 739 59 742 61
rect 744 59 747 61
rect 739 57 747 59
rect 749 65 754 68
rect 749 61 757 65
rect 749 59 752 61
rect 754 59 757 61
rect 749 57 757 59
rect 739 52 744 57
rect 752 54 757 57
rect 759 63 766 65
rect 782 67 784 69
rect 786 67 788 69
rect 782 64 788 67
rect 759 61 762 63
rect 764 61 766 63
rect 759 54 766 61
rect 772 60 777 64
rect 770 58 777 60
rect 770 56 772 58
rect 774 56 777 58
rect 770 54 777 56
rect 779 61 788 64
rect 779 54 790 61
rect 792 58 799 61
rect 792 56 795 58
rect 797 56 799 58
rect 792 54 799 56
<< pdif >>
rect 9 320 14 327
rect 7 318 14 320
rect 7 316 9 318
rect 11 316 14 318
rect 7 314 14 316
rect 16 314 25 327
rect 18 310 25 314
rect 18 308 20 310
rect 22 308 25 310
rect 18 305 25 308
rect 27 318 35 327
rect 27 316 30 318
rect 32 316 35 318
rect 27 305 35 316
rect 37 325 45 327
rect 37 323 40 325
rect 42 323 45 325
rect 37 318 45 323
rect 37 316 40 318
rect 42 316 45 318
rect 37 311 45 316
rect 37 309 40 311
rect 42 309 45 311
rect 37 305 45 309
rect 47 325 59 327
rect 47 323 54 325
rect 56 323 59 325
rect 47 305 59 323
rect 61 317 66 327
rect 70 325 77 327
rect 70 323 72 325
rect 74 323 77 325
rect 70 321 77 323
rect 61 309 68 317
rect 72 314 77 321
rect 79 319 88 327
rect 109 320 114 327
rect 79 314 90 319
rect 81 309 90 314
rect 92 317 99 319
rect 92 315 95 317
rect 97 315 99 317
rect 92 313 99 315
rect 107 318 114 320
rect 107 316 109 318
rect 111 316 114 318
rect 107 314 114 316
rect 116 314 125 327
rect 92 309 97 313
rect 118 310 125 314
rect 61 307 64 309
rect 66 307 68 309
rect 61 305 68 307
rect 81 307 83 309
rect 85 307 88 309
rect 81 305 88 307
rect 118 308 120 310
rect 122 308 125 310
rect 118 305 125 308
rect 127 318 135 327
rect 127 316 130 318
rect 132 316 135 318
rect 127 305 135 316
rect 137 325 145 327
rect 137 323 140 325
rect 142 323 145 325
rect 137 318 145 323
rect 137 316 140 318
rect 142 316 145 318
rect 137 311 145 316
rect 137 309 140 311
rect 142 309 145 311
rect 137 305 145 309
rect 147 325 159 327
rect 147 323 154 325
rect 156 323 159 325
rect 147 305 159 323
rect 161 317 166 327
rect 170 325 177 327
rect 170 323 172 325
rect 174 323 177 325
rect 170 321 177 323
rect 161 309 168 317
rect 172 314 177 321
rect 179 319 188 327
rect 209 320 214 327
rect 179 314 190 319
rect 181 309 190 314
rect 192 317 199 319
rect 192 315 195 317
rect 197 315 199 317
rect 192 313 199 315
rect 207 318 214 320
rect 207 316 209 318
rect 211 316 214 318
rect 207 314 214 316
rect 216 314 225 327
rect 192 309 197 313
rect 218 310 225 314
rect 161 307 164 309
rect 166 307 168 309
rect 161 305 168 307
rect 181 307 183 309
rect 185 307 188 309
rect 181 305 188 307
rect 218 308 220 310
rect 222 308 225 310
rect 218 305 225 308
rect 227 318 235 327
rect 227 316 230 318
rect 232 316 235 318
rect 227 305 235 316
rect 237 325 245 327
rect 237 323 240 325
rect 242 323 245 325
rect 237 318 245 323
rect 237 316 240 318
rect 242 316 245 318
rect 237 311 245 316
rect 237 309 240 311
rect 242 309 245 311
rect 237 305 245 309
rect 247 325 259 327
rect 247 323 254 325
rect 256 323 259 325
rect 247 305 259 323
rect 261 317 266 327
rect 270 325 277 327
rect 270 323 272 325
rect 274 323 277 325
rect 270 321 277 323
rect 261 309 268 317
rect 272 314 277 321
rect 279 319 288 327
rect 309 320 314 327
rect 279 314 290 319
rect 281 309 290 314
rect 292 317 299 319
rect 292 315 295 317
rect 297 315 299 317
rect 292 313 299 315
rect 307 318 314 320
rect 307 316 309 318
rect 311 316 314 318
rect 307 314 314 316
rect 316 314 325 327
rect 292 309 297 313
rect 318 310 325 314
rect 261 307 264 309
rect 266 307 268 309
rect 261 305 268 307
rect 281 307 283 309
rect 285 307 288 309
rect 281 305 288 307
rect 318 308 320 310
rect 322 308 325 310
rect 318 305 325 308
rect 327 318 335 327
rect 327 316 330 318
rect 332 316 335 318
rect 327 305 335 316
rect 337 318 345 327
rect 337 316 340 318
rect 342 316 345 318
rect 337 311 345 316
rect 337 309 340 311
rect 342 309 345 311
rect 337 305 345 309
rect 347 325 359 327
rect 347 323 354 325
rect 356 323 359 325
rect 347 305 359 323
rect 361 317 366 327
rect 370 325 377 327
rect 370 323 372 325
rect 374 323 377 325
rect 370 321 377 323
rect 361 309 368 317
rect 372 314 377 321
rect 379 319 388 327
rect 409 320 414 327
rect 379 314 390 319
rect 381 309 390 314
rect 392 317 399 319
rect 392 315 395 317
rect 397 315 399 317
rect 392 313 399 315
rect 407 318 414 320
rect 407 316 409 318
rect 411 316 414 318
rect 407 314 414 316
rect 416 314 425 327
rect 392 309 397 313
rect 418 310 425 314
rect 361 307 364 309
rect 366 307 368 309
rect 361 305 368 307
rect 381 307 383 309
rect 385 307 388 309
rect 381 305 388 307
rect 418 308 420 310
rect 422 308 425 310
rect 418 305 425 308
rect 427 318 435 327
rect 427 316 430 318
rect 432 316 435 318
rect 427 305 435 316
rect 437 325 445 327
rect 437 323 440 325
rect 442 323 445 325
rect 437 318 445 323
rect 437 316 440 318
rect 442 316 445 318
rect 437 311 445 316
rect 437 309 440 311
rect 442 309 445 311
rect 437 305 445 309
rect 447 325 459 327
rect 447 323 454 325
rect 456 323 459 325
rect 447 305 459 323
rect 461 317 466 327
rect 470 325 477 327
rect 470 323 472 325
rect 474 323 477 325
rect 470 321 477 323
rect 461 309 468 317
rect 472 314 477 321
rect 479 319 488 327
rect 509 320 514 327
rect 479 314 490 319
rect 481 309 490 314
rect 492 317 499 319
rect 492 315 495 317
rect 497 315 499 317
rect 492 313 499 315
rect 507 318 514 320
rect 507 316 509 318
rect 511 316 514 318
rect 507 314 514 316
rect 516 314 525 327
rect 492 309 497 313
rect 518 310 525 314
rect 461 307 464 309
rect 466 307 468 309
rect 461 305 468 307
rect 481 307 483 309
rect 485 307 488 309
rect 481 305 488 307
rect 518 308 520 310
rect 522 308 525 310
rect 518 305 525 308
rect 527 318 535 327
rect 527 316 530 318
rect 532 316 535 318
rect 527 305 535 316
rect 537 325 545 327
rect 537 323 540 325
rect 542 323 545 325
rect 537 318 545 323
rect 537 316 540 318
rect 542 316 545 318
rect 537 311 545 316
rect 537 309 540 311
rect 542 309 545 311
rect 537 305 545 309
rect 547 325 559 327
rect 547 323 554 325
rect 556 323 559 325
rect 547 305 559 323
rect 561 317 566 327
rect 570 325 577 327
rect 570 323 572 325
rect 574 323 577 325
rect 570 321 577 323
rect 561 309 568 317
rect 572 314 577 321
rect 579 319 588 327
rect 609 320 614 327
rect 579 314 590 319
rect 581 309 590 314
rect 592 317 599 319
rect 592 315 595 317
rect 597 315 599 317
rect 592 313 599 315
rect 607 318 614 320
rect 607 316 609 318
rect 611 316 614 318
rect 607 314 614 316
rect 616 314 625 327
rect 592 309 597 313
rect 618 310 625 314
rect 561 307 564 309
rect 566 307 568 309
rect 561 305 568 307
rect 581 307 583 309
rect 585 307 588 309
rect 581 305 588 307
rect 618 308 620 310
rect 622 308 625 310
rect 618 305 625 308
rect 627 318 635 327
rect 627 316 630 318
rect 632 316 635 318
rect 627 305 635 316
rect 637 325 645 327
rect 637 323 640 325
rect 642 323 645 325
rect 637 318 645 323
rect 637 316 640 318
rect 642 316 645 318
rect 637 311 645 316
rect 637 309 640 311
rect 642 309 645 311
rect 637 305 645 309
rect 647 325 659 327
rect 647 323 654 325
rect 656 323 659 325
rect 647 305 659 323
rect 661 317 666 327
rect 670 325 677 327
rect 670 323 672 325
rect 674 323 677 325
rect 670 321 677 323
rect 661 309 668 317
rect 672 314 677 321
rect 679 319 688 327
rect 709 320 714 327
rect 679 314 690 319
rect 681 309 690 314
rect 692 317 699 319
rect 692 315 695 317
rect 697 315 699 317
rect 692 313 699 315
rect 707 318 714 320
rect 707 316 709 318
rect 711 316 714 318
rect 707 314 714 316
rect 716 314 725 327
rect 692 309 697 313
rect 718 310 725 314
rect 661 307 664 309
rect 666 307 668 309
rect 661 305 668 307
rect 681 307 683 309
rect 685 307 688 309
rect 681 305 688 307
rect 718 308 720 310
rect 722 308 725 310
rect 718 305 725 308
rect 727 318 735 327
rect 727 316 730 318
rect 732 316 735 318
rect 727 305 735 316
rect 737 325 745 327
rect 737 323 740 325
rect 742 323 745 325
rect 737 318 745 323
rect 737 316 740 318
rect 742 316 745 318
rect 737 311 745 316
rect 737 309 740 311
rect 742 309 745 311
rect 737 305 745 309
rect 747 325 759 327
rect 747 323 754 325
rect 756 323 759 325
rect 747 305 759 323
rect 761 317 766 327
rect 770 325 777 327
rect 770 323 772 325
rect 774 323 777 325
rect 770 321 777 323
rect 761 309 768 317
rect 772 314 777 321
rect 779 319 788 327
rect 779 314 790 319
rect 781 309 790 314
rect 792 317 799 319
rect 792 315 795 317
rect 797 315 799 317
rect 792 313 799 315
rect 792 309 797 313
rect 761 307 764 309
rect 766 307 768 309
rect 761 305 768 307
rect 781 307 783 309
rect 785 307 788 309
rect 781 305 788 307
rect 18 279 25 281
rect 18 277 21 279
rect 23 277 25 279
rect 38 279 45 281
rect 38 277 40 279
rect 42 277 45 279
rect 9 273 14 277
rect 7 271 14 273
rect 7 269 9 271
rect 11 269 14 271
rect 7 267 14 269
rect 16 272 25 277
rect 16 267 27 272
rect 18 259 27 267
rect 29 265 34 272
rect 38 269 45 277
rect 29 263 36 265
rect 29 261 32 263
rect 34 261 36 263
rect 29 259 36 261
rect 40 259 45 269
rect 47 263 59 281
rect 47 261 50 263
rect 52 261 59 263
rect 47 259 59 261
rect 61 277 69 281
rect 61 275 64 277
rect 66 275 69 277
rect 61 270 69 275
rect 61 268 64 270
rect 66 268 69 270
rect 61 263 69 268
rect 61 261 64 263
rect 66 261 69 263
rect 61 259 69 261
rect 71 270 79 281
rect 71 268 74 270
rect 76 268 79 270
rect 71 259 79 268
rect 81 278 88 281
rect 81 276 84 278
rect 86 276 88 278
rect 118 279 125 281
rect 118 277 121 279
rect 123 277 125 279
rect 138 279 145 281
rect 138 277 140 279
rect 142 277 145 279
rect 81 272 88 276
rect 109 273 114 277
rect 81 259 90 272
rect 92 270 99 272
rect 92 268 95 270
rect 97 268 99 270
rect 92 266 99 268
rect 107 271 114 273
rect 107 269 109 271
rect 111 269 114 271
rect 107 267 114 269
rect 116 272 125 277
rect 116 267 127 272
rect 92 259 97 266
rect 118 259 127 267
rect 129 265 134 272
rect 138 269 145 277
rect 129 263 136 265
rect 129 261 132 263
rect 134 261 136 263
rect 129 259 136 261
rect 140 259 145 269
rect 147 263 159 281
rect 147 261 150 263
rect 152 261 159 263
rect 147 259 159 261
rect 161 277 169 281
rect 161 275 164 277
rect 166 275 169 277
rect 161 270 169 275
rect 161 268 164 270
rect 166 268 169 270
rect 161 263 169 268
rect 161 261 164 263
rect 166 261 169 263
rect 161 259 169 261
rect 171 270 179 281
rect 171 268 174 270
rect 176 268 179 270
rect 171 259 179 268
rect 181 278 188 281
rect 181 276 184 278
rect 186 276 188 278
rect 218 279 225 281
rect 218 277 221 279
rect 223 277 225 279
rect 238 279 245 281
rect 238 277 240 279
rect 242 277 245 279
rect 181 272 188 276
rect 209 273 214 277
rect 181 259 190 272
rect 192 270 199 272
rect 192 268 195 270
rect 197 268 199 270
rect 192 266 199 268
rect 207 271 214 273
rect 207 269 209 271
rect 211 269 214 271
rect 207 267 214 269
rect 216 272 225 277
rect 216 267 227 272
rect 192 259 197 266
rect 218 259 227 267
rect 229 265 234 272
rect 238 269 245 277
rect 229 263 236 265
rect 229 261 232 263
rect 234 261 236 263
rect 229 259 236 261
rect 240 259 245 269
rect 247 263 259 281
rect 247 261 250 263
rect 252 261 259 263
rect 247 259 259 261
rect 261 277 269 281
rect 261 275 264 277
rect 266 275 269 277
rect 261 270 269 275
rect 261 268 264 270
rect 266 268 269 270
rect 261 263 269 268
rect 261 261 264 263
rect 266 261 269 263
rect 261 259 269 261
rect 271 270 279 281
rect 271 268 274 270
rect 276 268 279 270
rect 271 259 279 268
rect 281 278 288 281
rect 281 276 284 278
rect 286 276 288 278
rect 318 279 325 281
rect 318 277 321 279
rect 323 277 325 279
rect 338 279 345 281
rect 338 277 340 279
rect 342 277 345 279
rect 281 273 288 276
rect 309 273 314 277
rect 281 259 290 273
rect 292 271 299 273
rect 292 269 295 271
rect 297 269 299 271
rect 292 266 299 269
rect 307 271 314 273
rect 307 269 309 271
rect 311 269 314 271
rect 307 267 314 269
rect 316 272 325 277
rect 316 267 327 272
rect 292 259 297 266
rect 318 259 327 267
rect 329 265 334 272
rect 338 269 345 277
rect 329 263 336 265
rect 329 261 332 263
rect 334 261 336 263
rect 329 259 336 261
rect 340 259 345 269
rect 347 263 359 281
rect 347 261 350 263
rect 352 261 359 263
rect 347 259 359 261
rect 361 277 369 281
rect 361 275 364 277
rect 366 275 369 277
rect 361 270 369 275
rect 361 268 364 270
rect 366 268 369 270
rect 361 263 369 268
rect 361 261 364 263
rect 366 261 369 263
rect 361 259 369 261
rect 371 270 379 281
rect 371 268 374 270
rect 376 268 379 270
rect 371 259 379 268
rect 381 278 388 281
rect 381 276 384 278
rect 386 276 388 278
rect 420 279 427 281
rect 420 277 423 279
rect 425 277 427 279
rect 440 279 447 281
rect 440 277 442 279
rect 444 277 447 279
rect 381 272 388 276
rect 411 273 416 277
rect 381 259 390 272
rect 392 270 399 272
rect 392 268 395 270
rect 397 268 399 270
rect 392 266 399 268
rect 409 271 416 273
rect 409 269 411 271
rect 413 269 416 271
rect 409 267 416 269
rect 418 272 427 277
rect 418 267 429 272
rect 392 259 397 266
rect 420 259 429 267
rect 431 265 436 272
rect 440 269 447 277
rect 431 263 438 265
rect 431 261 434 263
rect 436 261 438 263
rect 431 259 438 261
rect 442 259 447 269
rect 449 263 461 281
rect 449 261 452 263
rect 454 261 461 263
rect 449 259 461 261
rect 463 277 471 281
rect 463 275 466 277
rect 468 275 471 277
rect 463 270 471 275
rect 463 268 466 270
rect 468 268 471 270
rect 463 263 471 268
rect 463 261 466 263
rect 468 261 471 263
rect 463 259 471 261
rect 473 270 481 281
rect 473 268 476 270
rect 478 268 481 270
rect 473 259 481 268
rect 483 278 490 281
rect 483 276 486 278
rect 488 276 490 278
rect 520 279 527 281
rect 520 277 523 279
rect 525 277 527 279
rect 540 279 547 281
rect 540 277 542 279
rect 544 277 547 279
rect 483 273 490 276
rect 511 273 516 277
rect 483 260 492 273
rect 494 271 501 273
rect 494 269 497 271
rect 499 269 501 271
rect 494 266 501 269
rect 509 271 516 273
rect 509 269 511 271
rect 513 269 516 271
rect 509 267 516 269
rect 518 272 527 277
rect 518 267 529 272
rect 494 260 499 266
rect 483 259 490 260
rect 520 259 529 267
rect 531 265 536 272
rect 540 269 547 277
rect 531 263 538 265
rect 531 261 534 263
rect 536 261 538 263
rect 531 259 538 261
rect 542 259 547 269
rect 549 263 561 281
rect 549 261 552 263
rect 554 261 561 263
rect 549 259 561 261
rect 563 277 571 281
rect 563 275 566 277
rect 568 275 571 277
rect 563 270 571 275
rect 563 268 566 270
rect 568 268 571 270
rect 563 263 571 268
rect 563 261 566 263
rect 568 261 571 263
rect 563 259 571 261
rect 573 270 581 281
rect 573 268 576 270
rect 578 268 581 270
rect 573 259 581 268
rect 583 278 590 281
rect 583 276 586 278
rect 588 276 590 278
rect 620 279 627 281
rect 620 277 623 279
rect 625 277 627 279
rect 640 279 647 281
rect 640 277 642 279
rect 644 277 647 279
rect 583 272 590 276
rect 611 273 616 277
rect 583 259 592 272
rect 594 270 601 272
rect 594 268 597 270
rect 599 268 601 270
rect 594 266 601 268
rect 609 271 616 273
rect 609 269 611 271
rect 613 269 616 271
rect 609 267 616 269
rect 618 272 627 277
rect 618 267 629 272
rect 594 259 599 266
rect 620 259 629 267
rect 631 265 636 272
rect 640 269 647 277
rect 631 263 638 265
rect 631 261 634 263
rect 636 261 638 263
rect 631 259 638 261
rect 642 259 647 269
rect 649 263 661 281
rect 649 261 652 263
rect 654 261 661 263
rect 649 259 661 261
rect 663 277 671 281
rect 663 275 666 277
rect 668 275 671 277
rect 663 270 671 275
rect 663 268 666 270
rect 668 268 671 270
rect 663 263 671 268
rect 663 261 666 263
rect 668 261 671 263
rect 663 259 671 261
rect 673 270 681 281
rect 673 268 676 270
rect 678 268 681 270
rect 673 259 681 268
rect 683 278 690 281
rect 683 276 686 278
rect 688 276 690 278
rect 720 279 727 281
rect 720 277 723 279
rect 725 277 727 279
rect 740 279 747 281
rect 740 277 742 279
rect 744 277 747 279
rect 683 273 690 276
rect 711 273 716 277
rect 683 260 692 273
rect 694 271 701 273
rect 694 269 697 271
rect 699 269 701 271
rect 694 266 701 269
rect 709 271 716 273
rect 709 269 711 271
rect 713 269 716 271
rect 709 267 716 269
rect 718 272 727 277
rect 718 267 729 272
rect 694 260 699 266
rect 683 259 690 260
rect 720 259 729 267
rect 731 265 736 272
rect 740 269 747 277
rect 731 263 738 265
rect 731 261 734 263
rect 736 261 738 263
rect 731 259 738 261
rect 742 259 747 269
rect 749 263 761 281
rect 749 261 752 263
rect 754 261 761 263
rect 749 259 761 261
rect 763 277 771 281
rect 763 275 766 277
rect 768 275 771 277
rect 763 270 771 275
rect 763 268 766 270
rect 768 268 771 270
rect 763 263 771 268
rect 763 261 766 263
rect 768 261 771 263
rect 763 259 771 261
rect 773 270 781 281
rect 773 268 776 270
rect 778 268 781 270
rect 773 259 781 268
rect 783 278 790 281
rect 783 276 786 278
rect 788 276 790 278
rect 783 272 790 276
rect 783 259 792 272
rect 794 270 801 272
rect 794 268 797 270
rect 799 268 801 270
rect 794 266 801 268
rect 794 259 799 266
rect 18 175 27 183
rect 7 173 14 175
rect 7 171 9 173
rect 11 171 14 173
rect 7 169 14 171
rect 9 165 14 169
rect 16 170 27 175
rect 29 181 36 183
rect 29 179 32 181
rect 34 179 36 181
rect 29 177 36 179
rect 29 170 34 177
rect 40 173 45 183
rect 16 165 25 170
rect 38 165 45 173
rect 18 163 21 165
rect 23 163 25 165
rect 18 161 25 163
rect 38 163 40 165
rect 42 163 45 165
rect 38 161 45 163
rect 47 181 59 183
rect 47 179 50 181
rect 52 179 59 181
rect 47 161 59 179
rect 61 181 69 183
rect 61 179 64 181
rect 66 179 69 181
rect 61 174 69 179
rect 61 172 64 174
rect 66 172 69 174
rect 61 167 69 172
rect 61 165 64 167
rect 66 165 69 167
rect 61 161 69 165
rect 71 174 79 183
rect 71 172 74 174
rect 76 172 79 174
rect 71 161 79 172
rect 81 170 90 183
rect 92 176 97 183
rect 92 174 99 176
rect 118 175 127 183
rect 92 172 95 174
rect 97 172 99 174
rect 92 170 99 172
rect 107 173 114 175
rect 107 171 109 173
rect 111 171 114 173
rect 81 166 88 170
rect 81 164 84 166
rect 86 164 88 166
rect 107 169 114 171
rect 109 165 114 169
rect 116 170 127 175
rect 129 181 136 183
rect 129 179 132 181
rect 134 179 136 181
rect 129 177 136 179
rect 129 170 134 177
rect 140 173 145 183
rect 116 165 125 170
rect 138 165 145 173
rect 81 161 88 164
rect 118 163 121 165
rect 123 163 125 165
rect 118 161 125 163
rect 138 163 140 165
rect 142 163 145 165
rect 138 161 145 163
rect 147 181 159 183
rect 147 179 150 181
rect 152 179 159 181
rect 147 161 159 179
rect 161 181 169 183
rect 161 179 164 181
rect 166 179 169 181
rect 161 174 169 179
rect 161 172 164 174
rect 166 172 169 174
rect 161 167 169 172
rect 161 165 164 167
rect 166 165 169 167
rect 161 161 169 165
rect 171 174 179 183
rect 171 172 174 174
rect 176 172 179 174
rect 171 161 179 172
rect 181 170 190 183
rect 192 176 197 183
rect 192 174 199 176
rect 218 175 227 183
rect 192 172 195 174
rect 197 172 199 174
rect 192 170 199 172
rect 207 173 214 175
rect 207 171 209 173
rect 211 171 214 173
rect 181 166 188 170
rect 181 164 184 166
rect 186 164 188 166
rect 207 169 214 171
rect 209 165 214 169
rect 216 170 227 175
rect 229 181 236 183
rect 229 179 232 181
rect 234 179 236 181
rect 229 177 236 179
rect 229 170 234 177
rect 240 173 245 183
rect 216 165 225 170
rect 238 165 245 173
rect 181 161 188 164
rect 218 163 221 165
rect 223 163 225 165
rect 218 161 225 163
rect 238 163 240 165
rect 242 163 245 165
rect 238 161 245 163
rect 247 181 259 183
rect 247 179 250 181
rect 252 179 259 181
rect 247 161 259 179
rect 261 181 269 183
rect 261 179 264 181
rect 266 179 269 181
rect 261 174 269 179
rect 261 172 264 174
rect 266 172 269 174
rect 261 167 269 172
rect 261 165 264 167
rect 266 165 269 167
rect 261 161 269 165
rect 271 174 279 183
rect 271 172 274 174
rect 276 172 279 174
rect 271 161 279 172
rect 281 170 290 183
rect 292 176 297 183
rect 292 174 299 176
rect 318 175 327 183
rect 292 172 295 174
rect 297 172 299 174
rect 292 170 299 172
rect 307 173 314 175
rect 307 171 309 173
rect 311 171 314 173
rect 281 166 288 170
rect 281 164 284 166
rect 286 164 288 166
rect 307 169 314 171
rect 309 165 314 169
rect 316 170 327 175
rect 329 181 336 183
rect 329 179 332 181
rect 334 179 336 181
rect 329 177 336 179
rect 329 170 334 177
rect 340 173 345 183
rect 316 165 325 170
rect 338 165 345 173
rect 281 161 288 164
rect 318 163 321 165
rect 323 163 325 165
rect 318 161 325 163
rect 338 163 340 165
rect 342 163 345 165
rect 338 161 345 163
rect 347 181 359 183
rect 347 179 350 181
rect 352 179 359 181
rect 347 161 359 179
rect 361 181 369 183
rect 361 179 364 181
rect 366 179 369 181
rect 361 174 369 179
rect 361 172 364 174
rect 366 172 369 174
rect 361 167 369 172
rect 361 165 364 167
rect 366 165 369 167
rect 361 161 369 165
rect 371 174 379 183
rect 371 172 374 174
rect 376 172 379 174
rect 371 161 379 172
rect 381 170 390 183
rect 392 176 397 183
rect 392 174 399 176
rect 420 175 429 183
rect 392 172 395 174
rect 397 172 399 174
rect 392 170 399 172
rect 409 173 416 175
rect 409 171 411 173
rect 413 171 416 173
rect 381 166 388 170
rect 381 164 384 166
rect 386 164 388 166
rect 409 169 416 171
rect 411 165 416 169
rect 418 170 429 175
rect 431 181 438 183
rect 431 179 434 181
rect 436 179 438 181
rect 431 177 438 179
rect 431 170 436 177
rect 442 173 447 183
rect 418 165 427 170
rect 440 165 447 173
rect 381 161 388 164
rect 420 163 423 165
rect 425 163 427 165
rect 420 161 427 163
rect 440 163 442 165
rect 444 163 447 165
rect 440 161 447 163
rect 449 181 461 183
rect 449 179 452 181
rect 454 179 461 181
rect 449 161 461 179
rect 463 181 471 183
rect 463 179 466 181
rect 468 179 471 181
rect 463 174 471 179
rect 463 172 466 174
rect 468 172 471 174
rect 463 167 471 172
rect 463 165 466 167
rect 468 165 471 167
rect 463 161 471 165
rect 473 174 481 183
rect 473 172 476 174
rect 478 172 481 174
rect 473 161 481 172
rect 483 170 492 183
rect 494 176 499 183
rect 494 174 501 176
rect 520 175 529 183
rect 494 172 497 174
rect 499 172 501 174
rect 494 170 501 172
rect 509 173 516 175
rect 509 171 511 173
rect 513 171 516 173
rect 483 166 490 170
rect 483 164 486 166
rect 488 164 490 166
rect 509 169 516 171
rect 511 165 516 169
rect 518 170 529 175
rect 531 181 538 183
rect 531 179 534 181
rect 536 179 538 181
rect 531 177 538 179
rect 531 170 536 177
rect 542 173 547 183
rect 518 165 527 170
rect 540 165 547 173
rect 483 161 490 164
rect 520 163 523 165
rect 525 163 527 165
rect 520 161 527 163
rect 540 163 542 165
rect 544 163 547 165
rect 540 161 547 163
rect 549 181 561 183
rect 549 179 552 181
rect 554 179 561 181
rect 549 161 561 179
rect 563 181 571 183
rect 563 179 566 181
rect 568 179 571 181
rect 563 174 571 179
rect 563 172 566 174
rect 568 172 571 174
rect 563 167 571 172
rect 563 165 566 167
rect 568 165 571 167
rect 563 161 571 165
rect 573 174 581 183
rect 573 172 576 174
rect 578 172 581 174
rect 573 161 581 172
rect 583 170 592 183
rect 594 176 599 183
rect 594 174 601 176
rect 620 175 629 183
rect 594 172 597 174
rect 599 172 601 174
rect 594 170 601 172
rect 609 173 616 175
rect 609 171 611 173
rect 613 171 616 173
rect 583 166 590 170
rect 583 164 586 166
rect 588 164 590 166
rect 609 169 616 171
rect 611 165 616 169
rect 618 170 629 175
rect 631 181 638 183
rect 631 179 634 181
rect 636 179 638 181
rect 631 177 638 179
rect 631 170 636 177
rect 642 173 647 183
rect 618 165 627 170
rect 640 165 647 173
rect 583 161 590 164
rect 620 163 623 165
rect 625 163 627 165
rect 620 161 627 163
rect 640 163 642 165
rect 644 163 647 165
rect 640 161 647 163
rect 649 181 661 183
rect 649 179 652 181
rect 654 179 661 181
rect 649 161 661 179
rect 663 181 671 183
rect 663 179 666 181
rect 668 179 671 181
rect 663 174 671 179
rect 663 172 666 174
rect 668 172 671 174
rect 663 167 671 172
rect 663 165 666 167
rect 668 165 671 167
rect 663 161 671 165
rect 673 174 681 183
rect 673 172 676 174
rect 678 172 681 174
rect 673 161 681 172
rect 683 170 692 183
rect 694 176 699 183
rect 694 174 701 176
rect 720 175 729 183
rect 694 172 697 174
rect 699 172 701 174
rect 694 170 701 172
rect 709 173 716 175
rect 709 171 711 173
rect 713 171 716 173
rect 683 166 690 170
rect 683 164 686 166
rect 688 164 690 166
rect 709 169 716 171
rect 711 165 716 169
rect 718 170 729 175
rect 731 181 738 183
rect 731 179 734 181
rect 736 179 738 181
rect 731 177 738 179
rect 731 170 736 177
rect 742 173 747 183
rect 718 165 727 170
rect 740 165 747 173
rect 683 161 690 164
rect 720 163 723 165
rect 725 163 727 165
rect 720 161 727 163
rect 740 163 742 165
rect 744 163 747 165
rect 740 161 747 163
rect 749 181 761 183
rect 749 179 752 181
rect 754 179 761 181
rect 749 161 761 179
rect 763 181 771 183
rect 763 179 766 181
rect 768 179 771 181
rect 763 174 771 179
rect 763 172 766 174
rect 768 172 771 174
rect 763 167 771 172
rect 763 165 766 167
rect 768 165 771 167
rect 763 161 771 165
rect 773 174 781 183
rect 773 172 776 174
rect 778 172 781 174
rect 773 161 781 172
rect 783 170 792 183
rect 794 176 799 183
rect 794 174 801 176
rect 794 172 797 174
rect 799 172 801 174
rect 794 170 801 172
rect 783 166 790 170
rect 783 164 786 166
rect 788 164 790 166
rect 783 161 790 164
rect 18 135 25 137
rect 18 133 21 135
rect 23 133 25 135
rect 38 135 45 137
rect 38 133 40 135
rect 42 133 45 135
rect 9 129 14 133
rect 7 127 14 129
rect 7 125 9 127
rect 11 125 14 127
rect 7 123 14 125
rect 16 128 25 133
rect 16 123 27 128
rect 18 115 27 123
rect 29 121 34 128
rect 38 125 45 133
rect 29 119 36 121
rect 29 117 32 119
rect 34 117 36 119
rect 29 115 36 117
rect 40 115 45 125
rect 47 119 59 137
rect 47 117 50 119
rect 52 117 59 119
rect 47 115 59 117
rect 61 133 69 137
rect 61 131 64 133
rect 66 131 69 133
rect 61 126 69 131
rect 61 124 64 126
rect 66 124 69 126
rect 61 119 69 124
rect 61 117 64 119
rect 66 117 69 119
rect 61 115 69 117
rect 71 126 79 137
rect 71 124 74 126
rect 76 124 79 126
rect 71 115 79 124
rect 81 134 88 137
rect 81 132 84 134
rect 86 132 88 134
rect 118 135 125 137
rect 118 133 121 135
rect 123 133 125 135
rect 138 135 145 137
rect 138 133 140 135
rect 142 133 145 135
rect 81 128 88 132
rect 109 129 114 133
rect 81 115 90 128
rect 92 126 99 128
rect 92 124 95 126
rect 97 124 99 126
rect 92 122 99 124
rect 107 127 114 129
rect 107 125 109 127
rect 111 125 114 127
rect 107 123 114 125
rect 116 128 125 133
rect 116 123 127 128
rect 92 115 97 122
rect 118 115 127 123
rect 129 121 134 128
rect 138 125 145 133
rect 129 119 136 121
rect 129 117 132 119
rect 134 117 136 119
rect 129 115 136 117
rect 140 115 145 125
rect 147 119 159 137
rect 147 117 150 119
rect 152 117 159 119
rect 147 115 159 117
rect 161 133 169 137
rect 161 131 164 133
rect 166 131 169 133
rect 161 126 169 131
rect 161 124 164 126
rect 166 124 169 126
rect 161 119 169 124
rect 161 117 164 119
rect 166 117 169 119
rect 161 115 169 117
rect 171 126 179 137
rect 171 124 174 126
rect 176 124 179 126
rect 171 115 179 124
rect 181 134 188 137
rect 181 132 184 134
rect 186 132 188 134
rect 218 135 225 137
rect 218 133 221 135
rect 223 133 225 135
rect 238 135 245 137
rect 238 133 240 135
rect 242 133 245 135
rect 181 128 188 132
rect 209 129 214 133
rect 181 115 190 128
rect 192 126 199 128
rect 192 124 195 126
rect 197 124 199 126
rect 192 122 199 124
rect 207 127 214 129
rect 207 125 209 127
rect 211 125 214 127
rect 207 123 214 125
rect 216 128 225 133
rect 216 123 227 128
rect 192 115 197 122
rect 218 115 227 123
rect 229 121 234 128
rect 238 125 245 133
rect 229 119 236 121
rect 229 117 232 119
rect 234 117 236 119
rect 229 115 236 117
rect 240 115 245 125
rect 247 119 259 137
rect 247 117 250 119
rect 252 117 259 119
rect 247 115 259 117
rect 261 133 269 137
rect 261 131 264 133
rect 266 131 269 133
rect 261 126 269 131
rect 261 124 264 126
rect 266 124 269 126
rect 261 119 269 124
rect 261 117 264 119
rect 266 117 269 119
rect 261 115 269 117
rect 271 126 279 137
rect 271 124 274 126
rect 276 124 279 126
rect 271 115 279 124
rect 281 134 288 137
rect 281 132 284 134
rect 286 132 288 134
rect 318 135 325 137
rect 318 133 321 135
rect 323 133 325 135
rect 338 135 345 137
rect 338 133 340 135
rect 342 133 345 135
rect 281 128 288 132
rect 309 129 314 133
rect 281 115 290 128
rect 292 126 299 128
rect 292 124 295 126
rect 297 124 299 126
rect 292 122 299 124
rect 307 127 314 129
rect 307 125 309 127
rect 311 125 314 127
rect 307 123 314 125
rect 316 128 325 133
rect 316 123 327 128
rect 292 115 297 122
rect 318 115 327 123
rect 329 121 334 128
rect 338 125 345 133
rect 329 119 336 121
rect 329 117 332 119
rect 334 117 336 119
rect 329 115 336 117
rect 340 115 345 125
rect 347 119 359 137
rect 347 117 350 119
rect 352 117 359 119
rect 347 115 359 117
rect 361 133 369 137
rect 361 131 364 133
rect 366 131 369 133
rect 361 126 369 131
rect 361 124 364 126
rect 366 124 369 126
rect 361 119 369 124
rect 361 117 364 119
rect 366 117 369 119
rect 361 115 369 117
rect 371 126 379 137
rect 371 124 374 126
rect 376 124 379 126
rect 371 115 379 124
rect 381 134 388 137
rect 381 132 384 134
rect 386 132 388 134
rect 420 135 427 137
rect 420 133 423 135
rect 425 133 427 135
rect 440 135 447 137
rect 440 133 442 135
rect 444 133 447 135
rect 381 128 388 132
rect 411 129 416 133
rect 381 115 390 128
rect 392 126 399 128
rect 392 124 395 126
rect 397 124 399 126
rect 392 122 399 124
rect 409 127 416 129
rect 409 125 411 127
rect 413 125 416 127
rect 409 123 416 125
rect 418 128 427 133
rect 418 123 429 128
rect 392 115 397 122
rect 420 115 429 123
rect 431 121 436 128
rect 440 125 447 133
rect 431 119 438 121
rect 431 117 434 119
rect 436 117 438 119
rect 431 115 438 117
rect 442 115 447 125
rect 449 119 461 137
rect 449 117 452 119
rect 454 117 461 119
rect 449 115 461 117
rect 463 133 471 137
rect 463 131 466 133
rect 468 131 471 133
rect 463 126 471 131
rect 463 124 466 126
rect 468 124 471 126
rect 463 119 471 124
rect 463 117 466 119
rect 468 117 471 119
rect 463 115 471 117
rect 473 126 481 137
rect 473 124 476 126
rect 478 124 481 126
rect 473 115 481 124
rect 483 134 490 137
rect 483 132 486 134
rect 488 132 490 134
rect 520 135 527 137
rect 520 133 523 135
rect 525 133 527 135
rect 540 135 547 137
rect 540 133 542 135
rect 544 133 547 135
rect 483 128 490 132
rect 511 129 516 133
rect 483 115 492 128
rect 494 126 501 128
rect 494 124 497 126
rect 499 124 501 126
rect 494 122 501 124
rect 509 127 516 129
rect 509 125 511 127
rect 513 125 516 127
rect 509 123 516 125
rect 518 128 527 133
rect 518 123 529 128
rect 494 115 499 122
rect 520 115 529 123
rect 531 121 536 128
rect 540 125 547 133
rect 531 119 538 121
rect 531 117 534 119
rect 536 117 538 119
rect 531 115 538 117
rect 542 115 547 125
rect 549 119 561 137
rect 549 117 552 119
rect 554 117 561 119
rect 549 115 561 117
rect 563 133 571 137
rect 563 131 566 133
rect 568 131 571 133
rect 563 126 571 131
rect 563 124 566 126
rect 568 124 571 126
rect 563 119 571 124
rect 563 117 566 119
rect 568 117 571 119
rect 563 115 571 117
rect 573 126 581 137
rect 573 124 576 126
rect 578 124 581 126
rect 573 115 581 124
rect 583 134 590 137
rect 583 132 586 134
rect 588 132 590 134
rect 620 135 627 137
rect 620 133 623 135
rect 625 133 627 135
rect 640 135 647 137
rect 640 133 642 135
rect 644 133 647 135
rect 583 128 590 132
rect 611 129 616 133
rect 583 115 592 128
rect 594 126 601 128
rect 594 124 597 126
rect 599 124 601 126
rect 594 122 601 124
rect 609 127 616 129
rect 609 125 611 127
rect 613 125 616 127
rect 609 123 616 125
rect 618 128 627 133
rect 618 123 629 128
rect 594 115 599 122
rect 620 115 629 123
rect 631 121 636 128
rect 640 125 647 133
rect 631 119 638 121
rect 631 117 634 119
rect 636 117 638 119
rect 631 115 638 117
rect 642 115 647 125
rect 649 119 661 137
rect 649 117 652 119
rect 654 117 661 119
rect 649 115 661 117
rect 663 133 671 137
rect 663 131 666 133
rect 668 131 671 133
rect 663 126 671 131
rect 663 124 666 126
rect 668 124 671 126
rect 663 119 671 124
rect 663 117 666 119
rect 668 117 671 119
rect 663 115 671 117
rect 673 126 681 137
rect 673 124 676 126
rect 678 124 681 126
rect 673 115 681 124
rect 683 134 690 137
rect 683 132 686 134
rect 688 132 690 134
rect 720 135 727 137
rect 720 133 723 135
rect 725 133 727 135
rect 740 135 747 137
rect 740 133 742 135
rect 744 133 747 135
rect 683 128 690 132
rect 711 129 716 133
rect 683 115 692 128
rect 694 126 701 128
rect 694 124 697 126
rect 699 124 701 126
rect 694 122 701 124
rect 709 127 716 129
rect 709 125 711 127
rect 713 125 716 127
rect 709 123 716 125
rect 718 128 727 133
rect 718 123 729 128
rect 694 115 699 122
rect 720 115 729 123
rect 731 121 736 128
rect 740 125 747 133
rect 731 119 738 121
rect 731 117 734 119
rect 736 117 738 119
rect 731 115 738 117
rect 742 115 747 125
rect 749 119 761 137
rect 749 117 752 119
rect 754 117 761 119
rect 749 115 761 117
rect 763 133 771 137
rect 763 131 766 133
rect 768 131 771 133
rect 763 126 771 131
rect 763 124 766 126
rect 768 124 771 126
rect 763 119 771 124
rect 763 117 766 119
rect 768 117 771 119
rect 763 115 771 117
rect 773 126 781 137
rect 773 124 776 126
rect 778 124 781 126
rect 773 115 781 124
rect 783 134 790 137
rect 783 132 786 134
rect 788 132 790 134
rect 783 128 790 132
rect 783 115 792 128
rect 794 126 801 128
rect 794 124 797 126
rect 799 124 801 126
rect 794 122 801 124
rect 794 115 799 122
rect 9 32 14 39
rect 7 30 14 32
rect 7 28 9 30
rect 11 28 14 30
rect 7 26 14 28
rect 16 26 25 39
rect 18 22 25 26
rect 18 20 20 22
rect 22 20 25 22
rect 18 17 25 20
rect 27 30 35 39
rect 27 28 30 30
rect 32 28 35 30
rect 27 17 35 28
rect 37 37 45 39
rect 37 35 40 37
rect 42 35 45 37
rect 37 30 45 35
rect 37 28 40 30
rect 42 28 45 30
rect 37 23 45 28
rect 37 21 40 23
rect 42 21 45 23
rect 37 17 45 21
rect 47 37 59 39
rect 47 35 54 37
rect 56 35 59 37
rect 47 17 59 35
rect 61 29 66 39
rect 70 37 77 39
rect 70 35 72 37
rect 74 35 77 37
rect 70 33 77 35
rect 61 21 68 29
rect 72 26 77 33
rect 79 31 88 39
rect 109 32 114 39
rect 79 26 90 31
rect 81 21 90 26
rect 92 29 99 31
rect 92 27 95 29
rect 97 27 99 29
rect 92 25 99 27
rect 107 30 114 32
rect 107 28 109 30
rect 111 28 114 30
rect 107 26 114 28
rect 116 26 125 39
rect 92 21 97 25
rect 118 22 125 26
rect 61 19 64 21
rect 66 19 68 21
rect 61 17 68 19
rect 81 19 83 21
rect 85 19 88 21
rect 81 17 88 19
rect 118 20 120 22
rect 122 20 125 22
rect 118 17 125 20
rect 127 30 135 39
rect 127 28 130 30
rect 132 28 135 30
rect 127 17 135 28
rect 137 37 145 39
rect 137 35 140 37
rect 142 35 145 37
rect 137 30 145 35
rect 137 28 140 30
rect 142 28 145 30
rect 137 23 145 28
rect 137 21 140 23
rect 142 21 145 23
rect 137 17 145 21
rect 147 37 159 39
rect 147 35 154 37
rect 156 35 159 37
rect 147 17 159 35
rect 161 29 166 39
rect 170 37 177 39
rect 170 35 172 37
rect 174 35 177 37
rect 170 33 177 35
rect 161 21 168 29
rect 172 26 177 33
rect 179 31 188 39
rect 209 32 214 39
rect 179 26 190 31
rect 181 21 190 26
rect 192 29 199 31
rect 192 27 195 29
rect 197 27 199 29
rect 192 25 199 27
rect 207 30 214 32
rect 207 28 209 30
rect 211 28 214 30
rect 207 26 214 28
rect 216 26 225 39
rect 192 21 197 25
rect 218 22 225 26
rect 161 19 164 21
rect 166 19 168 21
rect 161 17 168 19
rect 181 19 183 21
rect 185 19 188 21
rect 181 17 188 19
rect 218 20 220 22
rect 222 20 225 22
rect 218 17 225 20
rect 227 30 235 39
rect 227 28 230 30
rect 232 28 235 30
rect 227 17 235 28
rect 237 37 245 39
rect 237 35 240 37
rect 242 35 245 37
rect 237 30 245 35
rect 237 28 240 30
rect 242 28 245 30
rect 237 23 245 28
rect 237 21 240 23
rect 242 21 245 23
rect 237 17 245 21
rect 247 37 259 39
rect 247 35 254 37
rect 256 35 259 37
rect 247 17 259 35
rect 261 29 266 39
rect 270 37 277 39
rect 270 35 272 37
rect 274 35 277 37
rect 270 33 277 35
rect 261 21 268 29
rect 272 26 277 33
rect 279 31 288 39
rect 309 32 314 39
rect 279 26 290 31
rect 281 21 290 26
rect 292 29 299 31
rect 292 27 295 29
rect 297 27 299 29
rect 292 25 299 27
rect 307 30 314 32
rect 307 28 309 30
rect 311 28 314 30
rect 307 26 314 28
rect 316 26 325 39
rect 292 21 297 25
rect 318 22 325 26
rect 261 19 264 21
rect 266 19 268 21
rect 261 17 268 19
rect 281 19 283 21
rect 285 19 288 21
rect 281 17 288 19
rect 318 20 320 22
rect 322 20 325 22
rect 318 17 325 20
rect 327 30 335 39
rect 327 28 330 30
rect 332 28 335 30
rect 327 17 335 28
rect 337 37 345 39
rect 337 35 340 37
rect 342 35 345 37
rect 337 30 345 35
rect 337 28 340 30
rect 342 28 345 30
rect 337 23 345 28
rect 337 21 340 23
rect 342 21 345 23
rect 337 17 345 21
rect 347 37 359 39
rect 347 35 354 37
rect 356 35 359 37
rect 347 17 359 35
rect 361 29 366 39
rect 370 37 377 39
rect 370 35 372 37
rect 374 35 377 37
rect 370 33 377 35
rect 361 21 368 29
rect 372 26 377 33
rect 379 31 388 39
rect 409 32 414 39
rect 379 26 390 31
rect 381 21 390 26
rect 392 29 399 31
rect 392 27 395 29
rect 397 27 399 29
rect 392 25 399 27
rect 407 30 414 32
rect 407 28 409 30
rect 411 28 414 30
rect 407 26 414 28
rect 416 26 425 39
rect 392 21 397 25
rect 418 22 425 26
rect 361 19 364 21
rect 366 19 368 21
rect 361 17 368 19
rect 381 19 383 21
rect 385 19 388 21
rect 381 17 388 19
rect 418 20 420 22
rect 422 20 425 22
rect 418 17 425 20
rect 427 30 435 39
rect 427 28 430 30
rect 432 28 435 30
rect 427 17 435 28
rect 437 37 445 39
rect 437 35 440 37
rect 442 35 445 37
rect 437 30 445 35
rect 437 28 440 30
rect 442 28 445 30
rect 437 23 445 28
rect 437 21 440 23
rect 442 21 445 23
rect 437 17 445 21
rect 447 37 459 39
rect 447 35 454 37
rect 456 35 459 37
rect 447 17 459 35
rect 461 29 466 39
rect 470 37 477 39
rect 470 35 472 37
rect 474 35 477 37
rect 470 33 477 35
rect 461 21 468 29
rect 472 26 477 33
rect 479 31 488 39
rect 509 32 514 39
rect 479 26 490 31
rect 481 21 490 26
rect 492 29 499 31
rect 492 27 495 29
rect 497 27 499 29
rect 492 25 499 27
rect 507 30 514 32
rect 507 28 509 30
rect 511 28 514 30
rect 507 26 514 28
rect 516 26 525 39
rect 492 21 497 25
rect 518 22 525 26
rect 461 19 464 21
rect 466 19 468 21
rect 461 17 468 19
rect 481 19 483 21
rect 485 19 488 21
rect 481 17 488 19
rect 518 20 520 22
rect 522 20 525 22
rect 518 17 525 20
rect 527 30 535 39
rect 527 28 530 30
rect 532 28 535 30
rect 527 17 535 28
rect 537 37 545 39
rect 537 35 540 37
rect 542 35 545 37
rect 537 30 545 35
rect 537 28 540 30
rect 542 28 545 30
rect 537 23 545 28
rect 537 21 540 23
rect 542 21 545 23
rect 537 17 545 21
rect 547 37 559 39
rect 547 35 554 37
rect 556 35 559 37
rect 547 17 559 35
rect 561 29 566 39
rect 570 37 577 39
rect 570 35 572 37
rect 574 35 577 37
rect 570 33 577 35
rect 561 21 568 29
rect 572 26 577 33
rect 579 31 588 39
rect 609 32 614 39
rect 579 26 590 31
rect 581 21 590 26
rect 592 29 599 31
rect 592 27 595 29
rect 597 27 599 29
rect 592 25 599 27
rect 607 30 614 32
rect 607 28 609 30
rect 611 28 614 30
rect 607 26 614 28
rect 616 26 625 39
rect 592 21 597 25
rect 618 22 625 26
rect 561 19 564 21
rect 566 19 568 21
rect 561 17 568 19
rect 581 19 583 21
rect 585 19 588 21
rect 581 17 588 19
rect 618 20 620 22
rect 622 20 625 22
rect 618 17 625 20
rect 627 30 635 39
rect 627 28 630 30
rect 632 28 635 30
rect 627 17 635 28
rect 637 37 645 39
rect 637 35 640 37
rect 642 35 645 37
rect 637 30 645 35
rect 637 28 640 30
rect 642 28 645 30
rect 637 23 645 28
rect 637 21 640 23
rect 642 21 645 23
rect 637 17 645 21
rect 647 37 659 39
rect 647 35 654 37
rect 656 35 659 37
rect 647 17 659 35
rect 661 29 666 39
rect 670 37 677 39
rect 670 35 672 37
rect 674 35 677 37
rect 670 33 677 35
rect 661 21 668 29
rect 672 26 677 33
rect 679 31 688 39
rect 709 32 714 39
rect 679 26 690 31
rect 681 21 690 26
rect 692 29 699 31
rect 692 27 695 29
rect 697 27 699 29
rect 692 25 699 27
rect 707 30 714 32
rect 707 28 709 30
rect 711 28 714 30
rect 707 26 714 28
rect 716 26 725 39
rect 692 21 697 25
rect 718 22 725 26
rect 661 19 664 21
rect 666 19 668 21
rect 661 17 668 19
rect 681 19 683 21
rect 685 19 688 21
rect 681 17 688 19
rect 718 20 720 22
rect 722 20 725 22
rect 718 17 725 20
rect 727 30 735 39
rect 727 28 730 30
rect 732 28 735 30
rect 727 17 735 28
rect 737 37 745 39
rect 737 35 740 37
rect 742 35 745 37
rect 737 30 745 35
rect 737 28 740 30
rect 742 28 745 30
rect 737 23 745 28
rect 737 21 740 23
rect 742 21 745 23
rect 737 17 745 21
rect 747 37 759 39
rect 747 35 754 37
rect 756 35 759 37
rect 747 17 759 35
rect 761 29 766 39
rect 770 37 777 39
rect 770 35 772 37
rect 774 35 777 37
rect 770 33 777 35
rect 761 21 768 29
rect 772 26 777 33
rect 779 31 788 39
rect 779 26 790 31
rect 781 21 790 26
rect 792 29 799 31
rect 792 27 795 29
rect 797 27 799 29
rect 792 25 799 27
rect 792 21 797 25
rect 761 19 764 21
rect 766 19 768 21
rect 761 17 768 19
rect 781 19 783 21
rect 785 19 788 21
rect 781 17 788 19
<< alu1 >>
rect 3 360 803 365
rect 3 358 10 360
rect 12 358 17 360
rect 19 358 110 360
rect 112 358 117 360
rect 119 358 210 360
rect 212 358 217 360
rect 219 358 310 360
rect 312 358 317 360
rect 319 358 410 360
rect 412 358 417 360
rect 419 358 510 360
rect 512 358 517 360
rect 519 358 610 360
rect 612 358 617 360
rect 619 358 710 360
rect 712 358 717 360
rect 719 358 803 360
rect 3 357 803 358
rect 79 351 83 357
rect 39 349 46 350
rect 39 347 42 349
rect 44 347 46 349
rect 39 346 46 347
rect 7 334 19 336
rect 7 332 14 334
rect 16 332 19 334
rect 7 330 19 332
rect 7 325 11 330
rect 7 323 8 325
rect 10 323 11 325
rect 7 322 11 323
rect 39 325 43 346
rect 39 323 40 325
rect 42 323 43 325
rect 39 318 43 323
rect 39 316 40 318
rect 42 316 43 318
rect 39 311 43 316
rect 79 342 83 347
rect 79 340 80 342
rect 82 340 83 342
rect 79 336 83 340
rect 76 335 83 336
rect 76 333 78 335
rect 80 333 83 335
rect 87 341 91 351
rect 139 349 146 350
rect 139 347 142 349
rect 144 347 146 349
rect 139 346 146 347
rect 179 350 183 351
rect 179 348 180 350
rect 182 348 183 350
rect 87 339 88 341
rect 90 339 91 341
rect 87 337 91 339
rect 87 335 88 337
rect 90 335 91 337
rect 87 333 91 335
rect 76 332 83 333
rect 79 328 83 332
rect 79 322 91 328
rect 107 334 119 336
rect 107 332 114 334
rect 116 332 119 334
rect 107 330 119 332
rect 107 326 111 330
rect 107 324 108 326
rect 110 324 111 326
rect 107 323 111 324
rect 107 318 111 319
rect 107 316 109 318
rect 107 315 111 316
rect 139 325 143 346
rect 139 323 140 325
rect 142 323 143 325
rect 139 322 143 323
rect 139 320 140 322
rect 142 320 143 322
rect 139 318 143 320
rect 139 316 140 318
rect 142 316 143 318
rect 139 311 143 316
rect 179 336 183 348
rect 176 335 183 336
rect 176 333 178 335
rect 180 333 183 335
rect 187 341 191 351
rect 239 349 246 350
rect 239 347 242 349
rect 244 347 246 349
rect 239 346 246 347
rect 279 349 283 350
rect 187 339 188 341
rect 190 339 191 341
rect 187 337 191 339
rect 187 335 188 337
rect 190 335 191 337
rect 187 333 191 335
rect 176 332 183 333
rect 179 328 183 332
rect 179 322 191 328
rect 207 334 219 336
rect 207 332 214 334
rect 216 332 219 334
rect 207 330 219 332
rect 207 325 211 330
rect 207 323 208 325
rect 210 323 211 325
rect 207 322 211 323
rect 239 329 243 346
rect 239 327 240 329
rect 242 327 243 329
rect 239 325 243 327
rect 239 323 240 325
rect 242 323 243 325
rect 239 318 243 323
rect 239 316 240 318
rect 242 316 243 318
rect 239 311 243 316
rect 279 347 280 349
rect 282 347 283 349
rect 279 336 283 347
rect 276 335 283 336
rect 276 333 278 335
rect 280 333 283 335
rect 287 341 291 351
rect 339 349 346 350
rect 339 347 342 349
rect 344 347 346 349
rect 339 346 346 347
rect 287 339 288 341
rect 290 339 291 341
rect 287 337 291 339
rect 287 335 288 337
rect 290 335 291 337
rect 287 333 291 335
rect 276 332 283 333
rect 279 328 283 332
rect 279 322 291 328
rect 307 334 319 336
rect 307 333 314 334
rect 307 331 308 333
rect 310 332 314 333
rect 316 332 319 334
rect 310 331 319 332
rect 307 330 319 331
rect 307 322 311 330
rect 339 325 343 346
rect 339 323 340 325
rect 342 323 343 325
rect 339 318 343 323
rect 339 316 340 318
rect 342 316 343 318
rect 339 311 343 316
rect 378 347 391 351
rect 387 341 391 347
rect 439 349 446 350
rect 439 347 442 349
rect 444 347 446 349
rect 439 346 446 347
rect 387 339 388 341
rect 390 339 391 341
rect 387 337 391 339
rect 376 335 383 336
rect 376 333 378 335
rect 380 333 383 335
rect 387 335 388 337
rect 390 335 391 337
rect 387 333 391 335
rect 376 332 383 333
rect 379 328 383 332
rect 379 325 391 328
rect 379 323 388 325
rect 390 323 391 325
rect 379 322 391 323
rect 407 334 419 336
rect 407 332 414 334
rect 416 332 419 334
rect 407 330 419 332
rect 407 325 411 330
rect 407 323 408 325
rect 410 323 411 325
rect 407 322 411 323
rect 439 325 443 346
rect 439 323 440 325
rect 442 323 443 325
rect 439 321 443 323
rect 439 319 440 321
rect 442 319 443 321
rect 439 318 443 319
rect 439 316 440 318
rect 442 316 443 318
rect 439 311 443 316
rect 478 347 491 351
rect 502 349 506 350
rect 487 341 491 347
rect 487 339 488 341
rect 490 339 491 341
rect 487 337 491 339
rect 476 335 483 336
rect 476 333 478 335
rect 480 333 483 335
rect 487 335 488 337
rect 490 335 491 337
rect 487 333 491 335
rect 476 332 483 333
rect 479 331 483 332
rect 479 329 480 331
rect 482 329 483 331
rect 479 328 483 329
rect 479 322 491 328
rect 502 347 503 349
rect 505 347 506 349
rect 502 336 506 347
rect 539 349 546 350
rect 539 347 542 349
rect 544 347 546 349
rect 539 346 546 347
rect 502 334 519 336
rect 502 332 514 334
rect 516 332 519 334
rect 507 330 519 332
rect 507 322 511 330
rect 539 333 543 346
rect 539 331 540 333
rect 542 331 543 333
rect 539 325 543 331
rect 539 323 540 325
rect 542 323 543 325
rect 539 318 543 323
rect 539 316 540 318
rect 542 316 543 318
rect 539 311 543 316
rect 578 347 591 351
rect 602 350 606 351
rect 602 348 603 350
rect 605 348 606 350
rect 587 341 591 347
rect 587 339 588 341
rect 590 339 591 341
rect 587 337 591 339
rect 576 335 583 336
rect 576 333 578 335
rect 580 333 583 335
rect 587 335 588 337
rect 590 335 591 337
rect 587 333 591 335
rect 576 332 583 333
rect 579 328 583 332
rect 579 325 591 328
rect 579 323 588 325
rect 590 323 591 325
rect 579 322 591 323
rect 602 336 606 348
rect 639 349 646 350
rect 639 347 642 349
rect 644 347 646 349
rect 639 346 646 347
rect 602 334 619 336
rect 602 332 614 334
rect 616 332 619 334
rect 607 330 619 332
rect 607 322 611 330
rect 639 333 643 346
rect 639 331 640 333
rect 642 331 643 333
rect 639 325 643 331
rect 639 323 640 325
rect 642 323 643 325
rect 639 318 643 323
rect 639 316 640 318
rect 642 316 643 318
rect 639 311 643 316
rect 678 347 691 351
rect 702 349 707 350
rect 687 341 691 347
rect 687 339 688 341
rect 690 339 691 341
rect 687 337 691 339
rect 676 335 683 336
rect 676 333 678 335
rect 680 333 683 335
rect 687 335 688 337
rect 690 335 691 337
rect 687 333 691 335
rect 676 332 683 333
rect 679 328 683 332
rect 679 325 691 328
rect 679 323 688 325
rect 690 323 691 325
rect 679 322 691 323
rect 702 347 704 349
rect 706 347 707 349
rect 702 336 707 347
rect 739 349 746 350
rect 739 347 742 349
rect 744 347 746 349
rect 739 346 746 347
rect 702 334 719 336
rect 702 332 714 334
rect 716 332 719 334
rect 707 330 719 332
rect 707 322 711 330
rect 739 325 743 346
rect 739 323 740 325
rect 742 323 743 325
rect 739 318 743 323
rect 739 316 740 318
rect 742 316 743 318
rect 739 311 743 316
rect 778 347 791 351
rect 787 341 791 347
rect 787 339 788 341
rect 790 339 791 341
rect 787 337 791 339
rect 776 335 783 336
rect 776 333 778 335
rect 780 333 783 335
rect 787 335 788 337
rect 790 335 791 337
rect 787 333 791 335
rect 776 332 783 333
rect 779 328 783 332
rect 779 325 791 328
rect 779 323 788 325
rect 790 323 791 325
rect 779 322 791 323
rect 30 310 40 311
rect 30 308 31 310
rect 33 309 40 310
rect 42 309 43 311
rect 33 308 43 309
rect 30 307 43 308
rect 130 309 140 311
rect 142 309 143 311
rect 130 307 143 309
rect 230 309 240 311
rect 242 309 243 311
rect 230 307 243 309
rect 330 309 340 311
rect 342 309 343 311
rect 330 307 343 309
rect 430 309 440 311
rect 442 309 443 311
rect 430 307 443 309
rect 530 309 540 311
rect 542 309 543 311
rect 530 307 543 309
rect 630 309 640 311
rect 642 309 643 311
rect 630 307 643 309
rect 730 310 740 311
rect 730 308 731 310
rect 733 309 740 310
rect 742 309 743 311
rect 733 308 743 309
rect 730 307 743 308
rect 3 300 803 301
rect 3 298 10 300
rect 12 298 110 300
rect 112 298 210 300
rect 212 298 310 300
rect 312 298 410 300
rect 412 298 510 300
rect 512 298 610 300
rect 612 298 710 300
rect 712 298 803 300
rect 3 293 803 298
rect 3 288 805 293
rect 3 286 94 288
rect 96 286 194 288
rect 196 286 294 288
rect 296 286 394 288
rect 396 286 496 288
rect 498 286 596 288
rect 598 286 696 288
rect 698 286 796 288
rect 798 286 805 288
rect 3 285 805 286
rect 63 277 76 279
rect 63 275 64 277
rect 66 275 76 277
rect 163 277 176 279
rect 163 275 164 277
rect 166 275 176 277
rect 263 277 276 279
rect 263 275 264 277
rect 266 275 276 277
rect 363 277 376 279
rect 363 275 364 277
rect 366 275 376 277
rect 465 277 478 279
rect 465 275 466 277
rect 468 275 478 277
rect 565 277 578 279
rect 565 275 566 277
rect 568 275 578 277
rect 665 277 678 279
rect 665 275 666 277
rect 668 275 678 277
rect 765 277 778 279
rect 765 275 766 277
rect 768 275 778 277
rect 15 258 27 264
rect 23 256 27 258
rect 23 254 24 256
rect 26 254 27 256
rect 23 253 30 254
rect 15 251 19 253
rect 15 249 16 251
rect 18 249 19 251
rect 23 251 26 253
rect 28 251 30 253
rect 23 250 30 251
rect 15 247 19 249
rect 15 245 16 247
rect 18 245 19 247
rect 15 239 19 245
rect 15 235 28 239
rect 63 270 67 275
rect 63 268 64 270
rect 66 268 67 270
rect 63 263 67 268
rect 63 261 64 263
rect 66 261 67 263
rect 63 240 67 261
rect 95 256 99 264
rect 87 254 99 256
rect 87 252 90 254
rect 92 252 104 254
rect 87 250 104 252
rect 60 239 68 240
rect 60 237 62 239
rect 64 237 65 239
rect 67 237 68 239
rect 60 236 68 237
rect 100 239 104 250
rect 100 237 101 239
rect 103 237 104 239
rect 115 264 119 265
rect 115 262 116 264
rect 118 262 127 264
rect 115 258 127 262
rect 123 254 127 258
rect 123 253 130 254
rect 115 251 119 253
rect 115 249 116 251
rect 118 249 119 251
rect 123 251 126 253
rect 128 251 130 253
rect 123 250 130 251
rect 115 247 119 249
rect 115 245 116 247
rect 118 245 119 247
rect 115 239 119 245
rect 100 236 104 237
rect 115 235 128 239
rect 163 270 167 275
rect 163 268 164 270
rect 166 268 167 270
rect 163 263 167 268
rect 163 261 164 263
rect 166 261 167 263
rect 163 240 167 261
rect 195 263 204 264
rect 195 261 201 263
rect 203 261 204 263
rect 195 260 204 261
rect 195 257 199 260
rect 192 256 199 257
rect 187 254 193 256
rect 195 254 199 256
rect 187 252 190 254
rect 192 252 199 254
rect 187 250 199 252
rect 215 258 227 264
rect 223 256 227 258
rect 223 254 224 256
rect 226 254 227 256
rect 223 253 230 254
rect 215 251 219 253
rect 215 249 216 251
rect 218 249 219 251
rect 223 251 226 253
rect 228 251 230 253
rect 223 250 230 251
rect 215 247 219 249
rect 215 245 216 247
rect 218 245 219 247
rect 160 239 168 240
rect 160 237 162 239
rect 164 237 165 239
rect 167 237 168 239
rect 160 236 168 237
rect 215 239 219 245
rect 215 235 228 239
rect 263 270 267 275
rect 263 268 264 270
rect 266 268 267 270
rect 263 263 267 268
rect 263 261 264 263
rect 266 261 267 263
rect 263 240 267 261
rect 295 264 304 265
rect 295 262 301 264
rect 303 262 304 264
rect 295 261 304 262
rect 295 256 299 261
rect 287 254 299 256
rect 287 252 290 254
rect 292 252 299 254
rect 287 250 299 252
rect 315 264 319 265
rect 315 262 316 264
rect 318 262 327 264
rect 315 258 327 262
rect 323 254 327 258
rect 323 253 330 254
rect 315 251 319 253
rect 315 249 316 251
rect 318 249 319 251
rect 323 251 326 253
rect 328 251 330 253
rect 323 250 330 251
rect 315 247 319 249
rect 315 245 316 247
rect 318 245 319 247
rect 260 239 268 240
rect 260 237 262 239
rect 264 237 265 239
rect 267 237 268 239
rect 260 236 268 237
rect 315 239 319 245
rect 315 235 328 239
rect 363 270 367 275
rect 363 268 364 270
rect 366 268 367 270
rect 363 263 367 268
rect 363 261 364 263
rect 366 261 367 263
rect 363 240 367 261
rect 395 257 399 264
rect 392 256 399 257
rect 387 254 393 256
rect 395 254 399 256
rect 387 252 390 254
rect 392 252 406 254
rect 387 250 406 252
rect 360 239 368 240
rect 360 237 362 239
rect 364 237 365 239
rect 367 237 368 239
rect 360 236 368 237
rect 402 239 406 250
rect 402 237 403 239
rect 405 237 406 239
rect 417 258 429 264
rect 425 256 429 258
rect 425 254 426 256
rect 428 254 429 256
rect 425 253 432 254
rect 417 251 421 253
rect 417 249 418 251
rect 420 249 421 251
rect 425 251 428 253
rect 430 251 432 253
rect 425 250 432 251
rect 417 247 421 249
rect 417 245 418 247
rect 420 245 421 247
rect 417 239 421 245
rect 402 235 406 237
rect 417 235 430 239
rect 465 270 469 275
rect 465 268 466 270
rect 468 268 469 270
rect 465 263 469 268
rect 465 261 466 263
rect 468 261 469 263
rect 465 240 469 261
rect 497 264 506 265
rect 497 262 503 264
rect 505 262 506 264
rect 497 261 506 262
rect 497 256 501 261
rect 489 254 501 256
rect 489 252 492 254
rect 494 252 501 254
rect 489 250 501 252
rect 517 264 521 265
rect 517 262 518 264
rect 520 262 529 264
rect 517 258 529 262
rect 525 254 529 258
rect 525 253 532 254
rect 517 251 521 253
rect 517 249 518 251
rect 520 249 521 251
rect 525 251 528 253
rect 530 251 532 253
rect 525 250 532 251
rect 517 247 521 249
rect 517 245 518 247
rect 520 245 521 247
rect 462 239 470 240
rect 462 237 464 239
rect 466 237 467 239
rect 469 237 470 239
rect 462 236 470 237
rect 517 239 521 245
rect 517 235 530 239
rect 565 270 569 275
rect 565 268 566 270
rect 568 268 569 270
rect 565 263 569 268
rect 565 261 566 263
rect 568 261 569 263
rect 565 240 569 261
rect 597 257 601 264
rect 594 256 601 257
rect 589 254 595 256
rect 597 254 601 256
rect 589 252 592 254
rect 594 252 601 254
rect 589 250 601 252
rect 617 258 629 264
rect 625 256 629 258
rect 625 254 626 256
rect 628 254 629 256
rect 625 253 632 254
rect 617 251 621 253
rect 617 249 618 251
rect 620 249 621 251
rect 625 251 628 253
rect 630 251 632 253
rect 625 250 632 251
rect 617 247 621 249
rect 617 245 618 247
rect 620 245 621 247
rect 562 239 570 240
rect 562 237 564 239
rect 566 237 567 239
rect 569 237 570 239
rect 562 236 570 237
rect 617 239 621 245
rect 617 235 630 239
rect 665 270 669 275
rect 665 268 666 270
rect 668 268 669 270
rect 665 263 669 268
rect 665 261 666 263
rect 668 261 669 263
rect 665 240 669 261
rect 697 264 706 265
rect 697 262 703 264
rect 705 262 706 264
rect 697 261 706 262
rect 697 256 701 261
rect 689 254 701 256
rect 689 252 692 254
rect 694 252 701 254
rect 689 250 701 252
rect 717 264 721 265
rect 717 262 718 264
rect 720 262 729 264
rect 717 258 729 262
rect 725 254 729 258
rect 725 253 732 254
rect 717 251 721 253
rect 717 249 718 251
rect 720 249 721 251
rect 725 251 728 253
rect 730 251 732 253
rect 725 250 732 251
rect 717 247 721 249
rect 717 245 718 247
rect 720 245 721 247
rect 662 239 670 240
rect 662 237 664 239
rect 666 237 667 239
rect 669 237 670 239
rect 662 236 670 237
rect 717 239 721 245
rect 717 235 730 239
rect 765 270 769 275
rect 765 268 766 270
rect 768 268 769 270
rect 765 263 769 268
rect 765 261 766 263
rect 768 261 769 263
rect 765 240 769 261
rect 797 257 801 264
rect 794 256 801 257
rect 789 254 795 256
rect 797 254 801 256
rect 789 252 792 254
rect 794 252 801 254
rect 789 250 801 252
rect 762 239 770 240
rect 762 237 764 239
rect 766 237 767 239
rect 769 237 770 239
rect 762 236 770 237
rect 3 228 805 229
rect 3 226 87 228
rect 89 226 94 228
rect 96 226 187 228
rect 189 226 194 228
rect 196 226 287 228
rect 289 226 294 228
rect 296 226 387 228
rect 389 226 394 228
rect 396 226 489 228
rect 491 226 496 228
rect 498 226 589 228
rect 591 226 596 228
rect 598 226 689 228
rect 691 226 696 228
rect 698 226 789 228
rect 791 226 796 228
rect 798 226 805 228
rect 3 216 805 226
rect 3 214 87 216
rect 89 214 94 216
rect 96 214 187 216
rect 189 214 194 216
rect 196 214 287 216
rect 289 214 294 216
rect 296 214 387 216
rect 389 214 394 216
rect 396 214 489 216
rect 491 214 496 216
rect 498 214 589 216
rect 591 214 596 216
rect 598 214 689 216
rect 691 214 696 216
rect 698 214 789 216
rect 791 214 796 216
rect 798 214 805 216
rect 3 213 805 214
rect 15 203 28 207
rect 15 197 19 203
rect 15 195 16 197
rect 18 195 19 197
rect 15 193 19 195
rect 15 191 16 193
rect 18 191 19 193
rect 15 189 19 191
rect 23 191 30 192
rect 23 189 26 191
rect 28 189 30 191
rect 23 188 30 189
rect 60 205 67 206
rect 60 203 62 205
rect 64 203 67 205
rect 60 202 67 203
rect 100 205 104 206
rect 100 203 101 205
rect 103 203 104 205
rect 23 184 27 188
rect 15 181 27 184
rect 15 179 16 181
rect 18 179 27 181
rect 15 178 27 179
rect 63 181 67 202
rect 63 179 64 181
rect 66 179 67 181
rect 63 174 67 179
rect 63 172 64 174
rect 66 172 67 174
rect 63 171 67 172
rect 100 192 104 203
rect 87 190 104 192
rect 87 188 90 190
rect 92 188 104 190
rect 115 203 128 207
rect 87 186 99 188
rect 95 178 99 186
rect 115 197 119 203
rect 115 195 116 197
rect 118 195 119 197
rect 115 193 119 195
rect 115 191 116 193
rect 118 191 119 193
rect 115 189 119 191
rect 123 192 130 193
rect 123 190 126 192
rect 128 190 130 192
rect 123 189 130 190
rect 123 187 124 189
rect 126 188 130 189
rect 160 205 167 206
rect 160 203 162 205
rect 164 203 167 205
rect 160 202 167 203
rect 126 187 127 188
rect 123 184 127 187
rect 115 178 127 184
rect 63 169 64 171
rect 66 169 67 171
rect 163 181 167 202
rect 163 179 164 181
rect 166 179 167 181
rect 163 174 167 179
rect 163 172 164 174
rect 166 172 167 174
rect 63 167 67 169
rect 163 167 167 172
rect 215 203 228 207
rect 187 190 199 192
rect 187 188 190 190
rect 192 188 199 190
rect 187 186 199 188
rect 195 181 199 186
rect 195 179 196 181
rect 198 179 199 181
rect 195 178 199 179
rect 215 197 219 203
rect 215 195 216 197
rect 218 195 219 197
rect 215 193 219 195
rect 215 191 216 193
rect 218 191 219 193
rect 215 189 219 191
rect 223 191 230 192
rect 223 189 226 191
rect 228 189 230 191
rect 223 188 230 189
rect 260 205 267 206
rect 260 203 262 205
rect 264 203 267 205
rect 260 202 267 203
rect 299 206 303 207
rect 299 204 300 206
rect 302 204 303 206
rect 223 184 227 188
rect 215 181 227 184
rect 215 179 216 181
rect 218 179 227 181
rect 215 178 227 179
rect 263 181 267 202
rect 263 179 264 181
rect 266 179 267 181
rect 263 174 267 179
rect 263 172 264 174
rect 266 172 267 174
rect 263 167 267 172
rect 299 192 303 204
rect 287 190 303 192
rect 287 188 290 190
rect 292 189 303 190
rect 292 188 296 189
rect 287 187 296 188
rect 298 187 303 189
rect 287 186 303 187
rect 315 203 328 207
rect 295 178 299 186
rect 315 197 319 203
rect 315 195 316 197
rect 318 195 319 197
rect 315 193 319 195
rect 315 191 316 193
rect 318 191 319 193
rect 315 189 319 191
rect 323 192 330 194
rect 323 190 326 192
rect 328 190 330 192
rect 323 189 330 190
rect 323 187 324 189
rect 326 188 330 189
rect 360 205 367 206
rect 360 203 362 205
rect 364 203 367 205
rect 360 202 367 203
rect 394 208 404 209
rect 394 206 395 208
rect 397 206 404 208
rect 394 205 404 206
rect 326 187 327 188
rect 323 184 327 187
rect 315 178 327 184
rect 363 181 367 202
rect 363 179 364 181
rect 366 179 367 181
rect 363 174 367 179
rect 363 172 364 174
rect 366 172 367 174
rect 363 167 367 172
rect 400 192 404 205
rect 387 190 404 192
rect 387 188 389 190
rect 391 188 404 190
rect 387 187 404 188
rect 417 203 430 207
rect 387 186 398 187
rect 394 181 398 186
rect 394 179 395 181
rect 397 179 398 181
rect 394 178 398 179
rect 417 197 421 203
rect 417 195 418 197
rect 420 195 421 197
rect 417 193 421 195
rect 417 191 418 193
rect 420 191 421 193
rect 417 189 421 191
rect 425 191 432 192
rect 425 189 428 191
rect 430 189 432 191
rect 425 188 432 189
rect 462 205 469 206
rect 462 203 464 205
rect 466 203 469 205
rect 462 202 469 203
rect 425 184 429 188
rect 417 181 429 184
rect 417 179 418 181
rect 420 179 429 181
rect 417 178 429 179
rect 465 181 469 202
rect 465 179 466 181
rect 468 179 469 181
rect 465 174 469 179
rect 465 172 466 174
rect 468 172 469 174
rect 465 167 469 172
rect 517 203 530 207
rect 489 190 501 192
rect 489 188 492 190
rect 494 189 501 190
rect 494 188 498 189
rect 489 187 498 188
rect 500 187 501 189
rect 489 186 501 187
rect 497 178 501 186
rect 517 197 521 203
rect 517 195 518 197
rect 520 195 521 197
rect 517 193 521 195
rect 517 191 518 193
rect 520 191 521 193
rect 517 189 521 191
rect 525 192 532 193
rect 525 190 528 192
rect 530 190 532 192
rect 525 189 532 190
rect 525 187 526 189
rect 528 188 532 189
rect 562 205 569 206
rect 562 203 564 205
rect 566 203 569 205
rect 562 202 569 203
rect 528 187 529 188
rect 525 184 529 187
rect 517 178 529 184
rect 565 181 569 202
rect 565 179 566 181
rect 568 179 569 181
rect 565 174 569 179
rect 565 172 566 174
rect 568 172 569 174
rect 565 167 569 172
rect 617 203 630 207
rect 589 190 601 192
rect 589 188 592 190
rect 594 188 601 190
rect 589 186 601 188
rect 597 181 601 186
rect 597 179 598 181
rect 600 179 601 181
rect 597 178 601 179
rect 617 197 621 203
rect 617 195 618 197
rect 620 195 621 197
rect 617 193 621 195
rect 617 191 618 193
rect 620 191 621 193
rect 617 189 621 191
rect 625 191 632 192
rect 625 189 628 191
rect 630 189 632 191
rect 625 188 632 189
rect 662 205 669 206
rect 662 203 664 205
rect 666 203 669 205
rect 662 202 669 203
rect 625 184 629 188
rect 617 181 629 184
rect 617 179 618 181
rect 620 179 629 181
rect 617 178 629 179
rect 665 181 669 202
rect 665 179 666 181
rect 668 179 669 181
rect 665 174 669 179
rect 665 172 666 174
rect 668 172 669 174
rect 665 167 669 172
rect 717 203 730 207
rect 689 190 701 192
rect 689 188 692 190
rect 694 189 701 190
rect 694 188 698 189
rect 689 187 698 188
rect 700 187 701 189
rect 689 186 701 187
rect 697 178 701 186
rect 717 197 721 203
rect 717 195 718 197
rect 720 195 721 197
rect 717 193 721 195
rect 717 191 718 193
rect 720 191 721 193
rect 717 189 721 191
rect 725 192 732 193
rect 725 190 728 192
rect 730 190 732 192
rect 725 189 732 190
rect 725 187 726 189
rect 728 188 732 189
rect 762 205 769 206
rect 762 203 764 205
rect 766 203 769 205
rect 762 202 769 203
rect 728 187 729 188
rect 725 184 729 187
rect 717 178 729 184
rect 765 181 769 202
rect 765 179 766 181
rect 768 179 769 181
rect 765 174 769 179
rect 765 172 766 174
rect 768 172 769 174
rect 765 167 769 172
rect 789 191 816 192
rect 789 190 813 191
rect 789 188 792 190
rect 794 189 813 190
rect 815 189 816 191
rect 794 188 816 189
rect 789 186 801 188
rect 797 182 801 186
rect 796 181 801 182
rect 796 179 797 181
rect 799 179 801 181
rect 796 178 801 179
rect 63 165 64 167
rect 66 165 76 167
rect 63 163 76 165
rect 163 165 164 167
rect 166 166 176 167
rect 166 165 173 166
rect 163 164 173 165
rect 175 164 176 166
rect 163 163 176 164
rect 263 165 264 167
rect 266 166 276 167
rect 266 165 273 166
rect 263 164 273 165
rect 275 164 276 166
rect 263 163 276 164
rect 363 165 364 167
rect 366 166 376 167
rect 366 165 373 166
rect 363 164 373 165
rect 375 164 376 166
rect 363 163 376 164
rect 465 165 466 167
rect 468 166 478 167
rect 468 165 475 166
rect 465 164 475 165
rect 477 164 478 166
rect 465 163 478 164
rect 565 165 566 167
rect 568 166 578 167
rect 568 165 575 166
rect 565 164 575 165
rect 577 164 578 166
rect 565 163 578 164
rect 665 165 666 167
rect 668 166 678 167
rect 668 165 675 166
rect 665 164 675 165
rect 677 164 678 166
rect 665 163 678 164
rect 765 165 766 167
rect 768 166 778 167
rect 768 165 775 166
rect 765 164 775 165
rect 777 164 778 166
rect 765 163 778 164
rect 3 156 805 157
rect 3 154 94 156
rect 96 154 194 156
rect 196 154 294 156
rect 296 154 394 156
rect 396 154 496 156
rect 498 154 596 156
rect 598 154 696 156
rect 698 154 796 156
rect 798 154 805 156
rect 3 144 805 154
rect 3 142 94 144
rect 96 142 194 144
rect 196 142 294 144
rect 296 142 394 144
rect 396 142 496 144
rect 498 142 596 144
rect 598 142 696 144
rect 698 142 796 144
rect 798 142 805 144
rect 3 141 805 142
rect 63 133 76 135
rect 63 131 64 133
rect 66 131 76 133
rect 163 133 176 135
rect 163 131 164 133
rect 166 131 176 133
rect 263 133 276 135
rect 263 131 264 133
rect 266 131 276 133
rect 363 133 376 135
rect 363 131 364 133
rect 366 131 376 133
rect 465 133 478 135
rect 465 131 466 133
rect 468 131 478 133
rect 565 133 578 135
rect 565 131 566 133
rect 568 131 578 133
rect 665 133 678 135
rect 665 131 666 133
rect 668 131 678 133
rect 765 133 778 135
rect 765 131 766 133
rect 768 131 778 133
rect 15 119 27 120
rect 15 117 16 119
rect 18 117 27 119
rect 15 114 27 117
rect 23 110 27 114
rect 23 109 30 110
rect 15 107 19 109
rect 15 105 16 107
rect 18 105 19 107
rect 23 107 26 109
rect 28 107 30 109
rect 23 106 30 107
rect 15 95 19 105
rect 15 94 28 95
rect 63 126 67 131
rect 63 124 64 126
rect 66 124 67 126
rect 63 119 67 124
rect 63 117 64 119
rect 66 117 67 119
rect 63 115 67 117
rect 63 113 64 115
rect 66 113 67 115
rect 63 96 67 113
rect 95 119 99 120
rect 95 117 96 119
rect 98 117 99 119
rect 95 112 99 117
rect 87 110 99 112
rect 87 108 90 110
rect 92 108 99 110
rect 87 106 99 108
rect 115 117 127 121
rect 123 112 127 117
rect 123 111 130 112
rect 123 109 124 111
rect 126 109 130 111
rect 115 107 119 109
rect 115 105 116 107
rect 118 105 119 107
rect 123 107 127 109
rect 129 107 130 109
rect 123 106 130 107
rect 15 92 25 94
rect 27 92 28 94
rect 15 91 28 92
rect 60 95 67 96
rect 60 93 62 95
rect 64 93 67 95
rect 60 92 67 93
rect 115 95 119 105
rect 115 94 128 95
rect 163 126 167 131
rect 263 130 267 131
rect 263 128 264 130
rect 266 128 267 130
rect 163 124 164 126
rect 166 124 167 126
rect 163 119 167 124
rect 163 117 164 119
rect 166 117 167 119
rect 163 103 167 117
rect 163 101 164 103
rect 166 101 167 103
rect 163 96 167 101
rect 195 119 203 120
rect 195 117 200 119
rect 202 117 203 119
rect 195 116 203 117
rect 195 112 199 116
rect 187 110 199 112
rect 187 108 190 110
rect 192 108 199 110
rect 187 106 199 108
rect 215 114 227 120
rect 223 110 227 114
rect 223 109 230 110
rect 215 107 219 109
rect 215 105 216 107
rect 218 105 219 107
rect 115 92 124 94
rect 126 92 128 94
rect 115 91 128 92
rect 160 95 167 96
rect 160 93 162 95
rect 164 93 167 95
rect 160 92 167 93
rect 215 95 219 105
rect 223 107 226 109
rect 228 107 230 109
rect 223 103 230 107
rect 223 101 224 103
rect 226 101 227 103
rect 223 100 227 101
rect 215 94 228 95
rect 263 126 267 128
rect 263 124 264 126
rect 266 124 267 126
rect 263 119 267 124
rect 263 117 264 119
rect 266 117 267 119
rect 263 96 267 117
rect 295 119 299 120
rect 295 117 296 119
rect 298 117 299 119
rect 295 112 299 117
rect 287 111 299 112
rect 287 110 296 111
rect 287 108 290 110
rect 292 109 296 110
rect 298 109 299 111
rect 292 108 299 109
rect 287 106 299 108
rect 315 119 327 120
rect 315 117 316 119
rect 318 117 327 119
rect 315 114 327 117
rect 323 110 327 114
rect 323 109 330 110
rect 315 107 319 109
rect 315 105 316 107
rect 318 105 319 107
rect 323 107 326 109
rect 328 107 330 109
rect 323 106 330 107
rect 215 92 224 94
rect 226 92 228 94
rect 215 91 228 92
rect 260 95 267 96
rect 260 93 262 95
rect 264 93 267 95
rect 260 92 267 93
rect 315 95 319 105
rect 315 94 328 95
rect 363 126 367 131
rect 363 124 364 126
rect 366 124 367 126
rect 363 119 367 124
rect 363 117 364 119
rect 366 117 367 119
rect 363 111 367 117
rect 363 109 364 111
rect 366 109 367 111
rect 363 96 367 109
rect 395 119 399 120
rect 395 117 396 119
rect 398 117 399 119
rect 395 112 399 117
rect 387 110 399 112
rect 387 108 390 110
rect 392 108 399 110
rect 387 106 399 108
rect 417 119 429 120
rect 417 117 418 119
rect 420 117 429 119
rect 417 114 429 117
rect 425 110 429 114
rect 425 109 432 110
rect 417 107 421 109
rect 417 105 418 107
rect 420 105 421 107
rect 425 107 428 109
rect 430 107 432 109
rect 425 106 432 107
rect 315 92 324 94
rect 326 92 328 94
rect 315 91 328 92
rect 360 95 367 96
rect 360 93 362 95
rect 364 93 367 95
rect 360 92 367 93
rect 417 95 421 105
rect 417 94 430 95
rect 465 126 469 131
rect 565 130 569 131
rect 565 128 566 130
rect 568 128 569 130
rect 665 130 669 131
rect 665 128 666 130
rect 668 128 669 130
rect 465 124 466 126
rect 468 124 469 126
rect 465 123 469 124
rect 465 121 466 123
rect 468 121 469 123
rect 465 119 469 121
rect 465 117 466 119
rect 468 117 469 119
rect 465 96 469 117
rect 497 119 501 120
rect 497 117 498 119
rect 500 117 501 119
rect 497 112 501 117
rect 489 110 501 112
rect 489 108 492 110
rect 494 108 501 110
rect 489 106 501 108
rect 517 114 529 120
rect 525 112 529 114
rect 525 110 526 112
rect 528 110 529 112
rect 525 109 532 110
rect 517 107 521 109
rect 517 105 518 107
rect 520 105 521 107
rect 525 107 528 109
rect 530 107 532 109
rect 525 106 532 107
rect 417 92 426 94
rect 428 92 430 94
rect 417 91 430 92
rect 462 95 469 96
rect 462 93 464 95
rect 466 93 469 95
rect 462 92 469 93
rect 517 95 521 105
rect 517 94 530 95
rect 565 126 569 128
rect 565 124 566 126
rect 568 124 569 126
rect 565 119 569 124
rect 565 117 566 119
rect 568 117 569 119
rect 565 96 569 117
rect 597 112 601 120
rect 589 110 601 112
rect 589 108 592 110
rect 594 108 605 110
rect 589 106 605 108
rect 601 103 605 106
rect 601 101 602 103
rect 604 101 605 103
rect 601 100 605 101
rect 617 120 621 121
rect 617 118 618 120
rect 620 118 629 120
rect 617 114 629 118
rect 625 110 629 114
rect 625 109 632 110
rect 617 107 621 109
rect 617 105 618 107
rect 620 105 621 107
rect 625 107 628 109
rect 630 107 632 109
rect 625 106 632 107
rect 517 92 527 94
rect 529 92 530 94
rect 517 91 530 92
rect 562 95 569 96
rect 562 93 564 95
rect 566 93 569 95
rect 562 92 569 93
rect 617 95 621 105
rect 617 94 630 95
rect 665 126 669 128
rect 665 124 666 126
rect 668 124 669 126
rect 665 119 669 124
rect 665 117 666 119
rect 668 117 669 119
rect 665 96 669 117
rect 697 119 706 120
rect 697 117 703 119
rect 705 117 706 119
rect 697 115 706 117
rect 697 113 701 115
rect 694 112 701 113
rect 689 110 695 112
rect 697 110 701 112
rect 689 108 692 110
rect 694 108 701 110
rect 689 106 701 108
rect 717 114 729 120
rect 725 110 729 114
rect 725 109 732 110
rect 717 107 721 109
rect 717 105 718 107
rect 720 105 721 107
rect 617 92 627 94
rect 629 92 630 94
rect 617 91 630 92
rect 662 95 669 96
rect 662 93 664 95
rect 666 93 669 95
rect 662 92 669 93
rect 717 95 721 105
rect 725 107 728 109
rect 730 107 732 109
rect 725 106 732 107
rect 725 104 726 106
rect 728 104 732 106
rect 725 103 732 104
rect 717 94 730 95
rect 765 126 769 131
rect 765 124 766 126
rect 768 124 769 126
rect 765 119 769 124
rect 765 117 766 119
rect 768 117 769 119
rect 765 98 769 117
rect 765 96 766 98
rect 768 96 769 98
rect 796 119 816 120
rect 796 117 797 119
rect 799 117 813 119
rect 815 117 816 119
rect 796 116 816 117
rect 797 112 801 116
rect 789 110 801 112
rect 789 108 792 110
rect 794 108 801 110
rect 789 106 801 108
rect 717 92 727 94
rect 729 92 730 94
rect 717 91 730 92
rect 762 95 769 96
rect 762 93 764 95
rect 766 93 769 95
rect 762 92 769 93
rect 3 84 805 85
rect 3 82 87 84
rect 89 82 94 84
rect 96 82 187 84
rect 189 82 194 84
rect 196 82 287 84
rect 289 82 294 84
rect 296 82 387 84
rect 389 82 394 84
rect 396 82 489 84
rect 491 82 496 84
rect 498 82 589 84
rect 591 82 596 84
rect 598 82 689 84
rect 691 82 696 84
rect 698 82 789 84
rect 791 82 796 84
rect 798 82 805 84
rect 3 77 805 82
rect 3 72 803 77
rect 3 70 10 72
rect 12 70 17 72
rect 19 70 110 72
rect 112 70 117 72
rect 119 70 210 72
rect 212 70 217 72
rect 219 70 310 72
rect 312 70 317 72
rect 319 70 410 72
rect 412 70 417 72
rect 419 70 510 72
rect 512 70 517 72
rect 519 70 610 72
rect 612 70 617 72
rect 619 70 710 72
rect 712 70 717 72
rect 719 70 803 72
rect 3 69 803 70
rect 79 63 83 69
rect 39 61 46 62
rect 39 59 42 61
rect 44 59 46 61
rect 39 58 46 59
rect 7 46 19 48
rect 7 44 14 46
rect 16 44 19 46
rect 7 42 19 44
rect 7 37 11 42
rect 7 35 8 37
rect 10 35 11 37
rect 7 34 11 35
rect 39 37 43 58
rect 39 35 40 37
rect 42 35 43 37
rect 39 30 43 35
rect 39 28 40 30
rect 42 28 43 30
rect 39 23 43 28
rect 79 54 83 59
rect 79 52 80 54
rect 82 52 83 54
rect 79 48 83 52
rect 76 47 83 48
rect 76 45 78 47
rect 80 45 83 47
rect 87 53 91 63
rect 139 61 146 62
rect 139 59 142 61
rect 144 59 146 61
rect 139 58 146 59
rect 179 62 183 63
rect 179 60 180 62
rect 182 60 183 62
rect 87 51 88 53
rect 90 51 91 53
rect 87 49 91 51
rect 87 47 88 49
rect 90 47 91 49
rect 87 45 91 47
rect 76 44 83 45
rect 79 40 83 44
rect 79 34 91 40
rect 107 46 119 48
rect 107 44 114 46
rect 116 44 119 46
rect 107 42 119 44
rect 107 38 111 42
rect 107 36 108 38
rect 110 36 111 38
rect 107 35 111 36
rect 107 30 111 31
rect 107 28 109 30
rect 107 27 111 28
rect 139 37 143 58
rect 139 35 140 37
rect 142 35 143 37
rect 139 30 143 35
rect 139 28 140 30
rect 142 28 143 30
rect 139 23 143 28
rect 179 48 183 60
rect 176 47 183 48
rect 176 45 178 47
rect 180 45 183 47
rect 187 53 191 63
rect 239 61 246 62
rect 239 59 242 61
rect 244 59 246 61
rect 239 58 246 59
rect 279 61 283 62
rect 187 51 188 53
rect 190 51 191 53
rect 187 49 191 51
rect 187 47 188 49
rect 190 47 191 49
rect 187 45 191 47
rect 176 44 183 45
rect 179 40 183 44
rect 179 34 191 40
rect 207 46 219 48
rect 207 44 214 46
rect 216 44 219 46
rect 207 42 219 44
rect 207 37 211 42
rect 207 35 208 37
rect 210 35 211 37
rect 207 34 211 35
rect 239 37 243 58
rect 239 35 240 37
rect 242 35 243 37
rect 239 30 243 35
rect 239 28 240 30
rect 242 28 243 30
rect 239 23 243 28
rect 279 59 280 61
rect 282 59 283 61
rect 279 48 283 59
rect 276 47 283 48
rect 276 45 278 47
rect 280 45 283 47
rect 287 53 291 63
rect 339 61 346 62
rect 339 59 342 61
rect 344 59 346 61
rect 339 58 346 59
rect 287 51 288 53
rect 290 51 291 53
rect 287 49 291 51
rect 287 47 288 49
rect 290 47 291 49
rect 287 45 291 47
rect 276 44 283 45
rect 279 40 283 44
rect 279 34 291 40
rect 307 46 319 48
rect 307 45 314 46
rect 307 43 308 45
rect 310 44 314 45
rect 316 44 319 46
rect 310 43 319 44
rect 307 42 319 43
rect 307 34 311 42
rect 339 37 343 58
rect 339 35 340 37
rect 342 35 343 37
rect 339 30 343 35
rect 339 28 340 30
rect 342 28 343 30
rect 339 23 343 28
rect 378 59 391 63
rect 387 53 391 59
rect 439 61 446 62
rect 439 59 442 61
rect 444 59 446 61
rect 439 58 446 59
rect 387 51 388 53
rect 390 51 391 53
rect 387 49 391 51
rect 376 47 383 48
rect 376 45 378 47
rect 380 45 383 47
rect 387 47 388 49
rect 390 47 391 49
rect 387 45 391 47
rect 376 44 383 45
rect 379 40 383 44
rect 379 37 391 40
rect 379 35 388 37
rect 390 35 391 37
rect 379 34 391 35
rect 407 46 419 48
rect 407 44 414 46
rect 416 44 419 46
rect 407 42 419 44
rect 407 37 411 42
rect 407 35 408 37
rect 410 35 411 37
rect 407 34 411 35
rect 439 37 443 58
rect 439 35 440 37
rect 442 35 443 37
rect 439 30 443 35
rect 439 28 440 30
rect 442 28 443 30
rect 439 23 443 28
rect 478 59 491 63
rect 502 61 506 62
rect 487 53 491 59
rect 487 51 488 53
rect 490 51 491 53
rect 487 49 491 51
rect 476 47 483 48
rect 476 45 478 47
rect 480 45 483 47
rect 487 47 488 49
rect 490 47 491 49
rect 487 45 491 47
rect 476 44 483 45
rect 479 43 483 44
rect 479 41 480 43
rect 482 41 483 43
rect 479 40 483 41
rect 479 34 491 40
rect 502 59 503 61
rect 505 59 506 61
rect 502 48 506 59
rect 539 61 546 62
rect 539 59 542 61
rect 544 59 546 61
rect 539 58 546 59
rect 502 46 519 48
rect 502 45 514 46
rect 502 44 508 45
rect 507 43 508 44
rect 510 44 514 45
rect 516 44 519 46
rect 510 43 519 44
rect 507 42 519 43
rect 507 34 511 42
rect 539 37 543 58
rect 539 35 540 37
rect 542 35 543 37
rect 539 30 543 35
rect 539 28 540 30
rect 542 28 543 30
rect 539 23 543 28
rect 578 59 591 63
rect 602 62 606 63
rect 602 60 603 62
rect 605 60 606 62
rect 587 53 591 59
rect 587 51 588 53
rect 590 51 591 53
rect 587 49 591 51
rect 576 47 583 48
rect 576 45 578 47
rect 580 45 583 47
rect 587 47 588 49
rect 590 47 591 49
rect 587 45 591 47
rect 576 44 583 45
rect 579 40 583 44
rect 579 37 591 40
rect 579 35 588 37
rect 590 35 591 37
rect 579 34 591 35
rect 602 48 606 60
rect 639 61 646 62
rect 639 59 642 61
rect 644 59 646 61
rect 639 58 646 59
rect 602 46 619 48
rect 602 44 614 46
rect 616 44 619 46
rect 607 42 619 44
rect 607 34 611 42
rect 639 37 643 58
rect 639 35 640 37
rect 642 35 643 37
rect 639 30 643 35
rect 639 28 640 30
rect 642 28 643 30
rect 639 23 643 28
rect 678 59 691 63
rect 702 61 707 62
rect 687 53 691 59
rect 687 51 688 53
rect 690 51 691 53
rect 687 49 691 51
rect 676 47 683 48
rect 676 45 678 47
rect 680 45 683 47
rect 687 47 688 49
rect 690 47 691 49
rect 687 45 691 47
rect 676 44 683 45
rect 679 40 683 44
rect 679 37 691 40
rect 679 35 688 37
rect 690 35 691 37
rect 679 34 691 35
rect 702 59 704 61
rect 706 59 707 61
rect 702 48 707 59
rect 739 61 746 62
rect 739 59 742 61
rect 744 59 746 61
rect 739 58 746 59
rect 702 46 719 48
rect 702 44 714 46
rect 716 44 719 46
rect 707 42 719 44
rect 707 34 711 42
rect 739 37 743 58
rect 739 35 740 37
rect 742 35 743 37
rect 739 30 743 35
rect 739 28 740 30
rect 742 28 743 30
rect 739 23 743 28
rect 778 59 791 63
rect 787 53 791 59
rect 787 51 788 53
rect 790 51 791 53
rect 787 49 791 51
rect 776 47 783 48
rect 776 45 778 47
rect 780 45 783 47
rect 787 47 788 49
rect 790 47 791 49
rect 787 45 791 47
rect 776 44 783 45
rect 779 40 783 44
rect 779 37 791 40
rect 779 35 788 37
rect 790 35 791 37
rect 779 34 791 35
rect 30 21 40 23
rect 42 21 43 23
rect 30 19 43 21
rect 130 21 140 23
rect 142 21 143 23
rect 130 19 143 21
rect 230 21 240 23
rect 242 21 243 23
rect 230 19 243 21
rect 330 21 340 23
rect 342 21 343 23
rect 330 19 343 21
rect 430 21 440 23
rect 442 21 443 23
rect 430 19 443 21
rect 530 21 540 23
rect 542 21 543 23
rect 530 19 543 21
rect 630 21 640 23
rect 642 21 643 23
rect 630 19 643 21
rect 730 21 740 23
rect 742 21 743 23
rect 730 19 743 21
rect 3 12 803 13
rect 3 10 10 12
rect 12 10 110 12
rect 112 10 210 12
rect 212 10 310 12
rect 312 10 410 12
rect 412 10 510 12
rect 512 10 610 12
rect 612 10 710 12
rect 712 10 803 12
rect 3 5 803 10
<< alu2 >>
rect 79 362 707 366
rect 79 342 83 362
rect 179 354 606 358
rect 179 350 183 354
rect 602 350 606 354
rect 179 348 180 350
rect 182 348 183 350
rect 179 347 183 348
rect 279 349 506 350
rect 279 347 280 349
rect 282 347 503 349
rect 505 347 506 349
rect 602 348 603 350
rect 605 348 606 350
rect 602 347 606 348
rect 703 349 707 362
rect 703 347 704 349
rect 706 347 707 349
rect 279 346 506 347
rect 703 346 707 347
rect 79 340 80 342
rect 82 340 83 342
rect 79 339 83 340
rect 87 341 824 342
rect 87 339 88 341
rect 90 339 188 341
rect 190 339 288 341
rect 290 339 388 341
rect 390 339 488 341
rect 490 339 588 341
rect 590 339 688 341
rect 690 339 788 341
rect 790 339 821 341
rect 823 339 824 341
rect 87 338 824 339
rect 307 333 483 334
rect 307 331 308 333
rect 310 331 483 333
rect 307 330 480 331
rect 239 329 303 330
rect 239 327 240 329
rect 242 327 300 329
rect 302 327 303 329
rect 479 329 480 330
rect 482 329 483 331
rect 539 333 602 334
rect 539 331 540 333
rect 542 331 599 333
rect 601 331 602 333
rect 539 330 602 331
rect 639 333 643 334
rect 639 331 640 333
rect 642 331 643 333
rect 479 328 483 329
rect 639 328 643 331
rect 107 326 111 327
rect 239 326 303 327
rect 639 326 640 328
rect 642 326 643 328
rect 7 325 11 326
rect 7 323 8 325
rect 10 323 11 325
rect 7 297 11 323
rect 107 324 108 326
rect 110 324 111 326
rect 30 310 34 311
rect 30 308 31 310
rect 33 308 34 310
rect 30 304 34 308
rect 30 302 31 304
rect 33 302 34 304
rect 30 301 34 302
rect 107 305 111 324
rect 207 325 211 326
rect 207 323 208 325
rect 210 323 211 325
rect 139 322 143 323
rect 139 320 140 322
rect 142 320 143 322
rect 139 315 143 320
rect 139 313 140 315
rect 142 313 143 315
rect 139 311 143 313
rect 207 313 211 323
rect 339 325 343 326
rect 339 323 340 325
rect 342 323 343 325
rect 339 320 343 323
rect 387 325 411 326
rect 387 323 388 325
rect 390 323 408 325
rect 410 323 411 325
rect 387 322 411 323
rect 439 325 443 326
rect 439 323 440 325
rect 442 323 443 325
rect 339 318 340 320
rect 342 318 343 320
rect 339 317 343 318
rect 439 321 443 323
rect 439 319 440 321
rect 442 319 443 321
rect 439 317 443 319
rect 587 325 591 326
rect 587 323 588 325
rect 590 323 591 325
rect 587 313 591 323
rect 639 319 643 326
rect 687 325 691 326
rect 687 323 688 325
rect 690 323 691 325
rect 207 309 591 313
rect 687 305 691 323
rect 787 325 791 326
rect 787 323 788 325
rect 790 323 791 325
rect 107 301 691 305
rect 730 310 734 311
rect 730 308 731 310
rect 733 308 734 310
rect 730 304 734 308
rect 730 302 731 304
rect 733 302 734 304
rect 730 301 734 302
rect 787 297 791 323
rect 7 293 791 297
rect 339 288 706 289
rect 339 286 340 288
rect 342 286 703 288
rect 705 286 706 288
rect 339 285 706 286
rect 115 277 806 281
rect 115 264 119 277
rect 115 262 116 264
rect 118 262 119 264
rect 115 261 119 262
rect 200 272 204 273
rect 200 270 201 272
rect 203 270 204 272
rect 200 263 204 270
rect 200 261 201 263
rect 203 261 204 263
rect 300 272 304 273
rect 300 270 301 272
rect 303 270 304 272
rect 300 264 304 270
rect 300 262 301 264
rect 303 262 304 264
rect 300 261 304 262
rect 315 264 319 277
rect 315 262 316 264
rect 318 262 319 264
rect 315 261 319 262
rect 497 264 506 265
rect 497 262 498 264
rect 500 262 503 264
rect 505 262 506 264
rect 497 261 506 262
rect 517 264 521 277
rect 517 262 518 264
rect 520 262 521 264
rect 517 261 521 262
rect 702 272 706 273
rect 702 270 703 272
rect 705 270 706 272
rect 702 264 706 270
rect 702 262 703 264
rect 705 262 706 264
rect 702 261 706 262
rect 717 264 721 277
rect 717 262 718 264
rect 720 262 721 264
rect 717 261 721 262
rect 200 260 204 261
rect 23 256 196 257
rect 23 254 24 256
rect 26 254 193 256
rect 195 254 196 256
rect 23 253 196 254
rect 223 256 396 257
rect 223 254 224 256
rect 226 254 393 256
rect 395 254 396 256
rect 223 253 396 254
rect 425 256 602 257
rect 425 254 426 256
rect 428 254 595 256
rect 597 254 599 256
rect 601 254 602 256
rect 425 253 602 254
rect 625 256 798 257
rect 625 254 626 256
rect 628 254 789 256
rect 791 254 795 256
rect 797 254 798 256
rect 625 253 798 254
rect 15 247 721 248
rect 15 245 16 247
rect 18 245 116 247
rect 118 245 216 247
rect 218 245 316 247
rect 318 245 418 247
rect 420 245 518 247
rect 520 245 618 247
rect 620 245 718 247
rect 720 245 721 247
rect 15 244 721 245
rect 63 239 68 240
rect 63 237 65 239
rect 67 237 68 239
rect 63 236 68 237
rect 100 239 104 240
rect 100 237 101 239
rect 103 237 104 239
rect 63 211 67 236
rect 100 235 104 237
rect 100 233 101 235
rect 103 233 104 235
rect 100 232 104 233
rect 164 239 168 240
rect 164 237 165 239
rect 167 237 168 239
rect 164 211 168 237
rect 264 239 268 240
rect 264 237 265 239
rect 267 237 268 239
rect 264 222 268 237
rect 264 220 265 222
rect 267 220 268 222
rect 264 219 268 220
rect 364 239 368 240
rect 364 237 365 239
rect 367 237 368 239
rect 63 207 104 211
rect 164 207 303 211
rect 100 205 104 207
rect 100 203 101 205
rect 103 203 104 205
rect 299 206 303 207
rect 299 204 300 206
rect 302 204 303 206
rect 364 209 368 237
rect 402 239 406 240
rect 402 237 403 239
rect 405 237 406 239
rect 402 232 406 237
rect 466 239 470 240
rect 466 237 467 239
rect 469 237 470 239
rect 466 235 470 237
rect 402 230 403 232
rect 405 230 406 232
rect 465 231 470 235
rect 402 223 406 230
rect 466 229 470 231
rect 566 239 570 240
rect 566 237 567 239
rect 569 237 570 239
rect 466 228 506 229
rect 466 226 503 228
rect 505 226 506 228
rect 466 225 506 226
rect 566 228 570 237
rect 566 226 567 228
rect 569 226 570 228
rect 566 225 570 226
rect 666 239 670 240
rect 666 237 667 239
rect 669 237 670 239
rect 666 220 670 237
rect 666 218 667 220
rect 669 218 670 220
rect 766 239 770 240
rect 766 237 767 239
rect 769 237 770 239
rect 766 221 770 237
rect 766 219 767 221
rect 769 219 770 221
rect 766 218 770 219
rect 666 217 670 218
rect 802 209 806 277
rect 364 208 398 209
rect 364 206 395 208
rect 397 206 398 208
rect 364 205 398 206
rect 402 208 806 209
rect 402 206 403 208
rect 405 206 806 208
rect 402 205 806 206
rect 299 203 303 204
rect 100 202 104 203
rect 15 197 721 198
rect 15 195 16 197
rect 18 195 116 197
rect 118 195 216 197
rect 218 195 316 197
rect 318 195 418 197
rect 420 195 518 197
rect 520 195 618 197
rect 620 195 718 197
rect 720 195 721 197
rect 15 194 721 195
rect 802 190 806 205
rect 812 221 816 222
rect 812 219 813 221
rect 815 219 816 221
rect 812 191 816 219
rect 123 189 299 190
rect 123 187 124 189
rect 126 187 296 189
rect 298 187 299 189
rect 123 186 299 187
rect 323 189 406 190
rect 323 187 324 189
rect 326 187 403 189
rect 405 187 406 189
rect 323 186 406 187
rect 497 189 506 190
rect 497 187 498 189
rect 500 187 503 189
rect 505 187 506 189
rect 497 186 506 187
rect 525 189 705 190
rect 525 187 526 189
rect 528 187 698 189
rect 700 187 702 189
rect 704 187 705 189
rect 525 186 705 187
rect 725 189 808 190
rect 725 187 726 189
rect 728 187 808 189
rect 812 189 813 191
rect 815 189 816 191
rect 812 188 816 189
rect 725 186 808 187
rect 15 181 206 182
rect 15 179 16 181
rect 18 179 196 181
rect 198 179 203 181
rect 205 179 206 181
rect 15 178 206 179
rect 215 181 398 182
rect 215 179 216 181
rect 218 179 395 181
rect 397 179 398 181
rect 215 178 398 179
rect 417 181 606 182
rect 417 179 418 181
rect 420 179 598 181
rect 600 179 603 181
rect 605 179 606 181
rect 417 178 606 179
rect 617 181 800 182
rect 617 179 618 181
rect 620 179 797 181
rect 799 179 800 181
rect 617 178 800 179
rect 63 171 67 172
rect 63 169 64 171
rect 66 169 67 171
rect 63 157 67 169
rect 172 166 203 167
rect 172 164 173 166
rect 175 164 200 166
rect 202 164 203 166
rect 172 163 203 164
rect 272 166 303 167
rect 272 164 273 166
rect 275 164 300 166
rect 302 164 303 166
rect 272 163 303 164
rect 372 166 406 167
rect 372 164 373 166
rect 375 164 403 166
rect 405 164 406 166
rect 372 163 406 164
rect 474 166 478 167
rect 474 164 475 166
rect 477 164 478 166
rect 474 157 478 164
rect 63 156 99 157
rect 63 154 96 156
rect 98 154 99 156
rect 63 153 99 154
rect 395 153 478 157
rect 574 166 578 167
rect 574 164 575 166
rect 577 164 578 166
rect 574 156 578 164
rect 674 166 706 167
rect 674 164 675 166
rect 677 164 703 166
rect 705 164 706 166
rect 674 163 706 164
rect 774 166 778 167
rect 774 164 775 166
rect 777 164 778 166
rect 574 154 575 156
rect 577 154 578 156
rect 574 153 578 154
rect 774 156 778 164
rect 774 154 775 156
rect 777 154 778 156
rect 774 153 778 154
rect 395 149 399 153
rect 15 145 399 149
rect 15 119 19 145
rect 199 140 319 141
rect 199 138 200 140
rect 202 138 319 140
rect 15 117 16 119
rect 18 117 19 119
rect 15 116 19 117
rect 95 137 99 138
rect 95 135 96 137
rect 98 135 99 137
rect 95 119 99 135
rect 95 117 96 119
rect 98 117 99 119
rect 95 116 99 117
rect 199 137 319 138
rect 199 119 203 137
rect 263 130 267 131
rect 263 128 264 130
rect 266 128 267 130
rect 263 123 267 128
rect 263 121 264 123
rect 266 121 267 123
rect 263 120 267 121
rect 199 117 200 119
rect 202 117 203 119
rect 199 116 203 117
rect 295 119 303 120
rect 295 117 296 119
rect 298 117 300 119
rect 302 117 303 119
rect 295 116 303 117
rect 315 119 319 137
rect 315 117 316 119
rect 318 117 319 119
rect 315 116 319 117
rect 395 119 399 145
rect 395 117 396 119
rect 398 117 399 119
rect 395 116 399 117
rect 417 145 800 149
rect 417 119 421 145
rect 497 140 621 141
rect 497 138 498 140
rect 500 138 621 140
rect 497 137 621 138
rect 417 117 418 119
rect 420 117 421 119
rect 417 116 421 117
rect 465 123 469 124
rect 465 121 466 123
rect 468 121 469 123
rect 63 115 67 116
rect 63 113 64 115
rect 66 113 67 115
rect 63 102 67 113
rect 123 111 299 112
rect 123 109 124 111
rect 126 109 296 111
rect 298 109 299 111
rect 123 108 299 109
rect 351 111 367 112
rect 351 109 352 111
rect 354 109 364 111
rect 366 109 367 111
rect 351 108 367 109
rect 465 111 469 121
rect 497 119 501 137
rect 497 117 498 119
rect 500 117 501 119
rect 497 116 501 117
rect 505 132 509 133
rect 505 130 506 132
rect 508 130 509 132
rect 465 109 466 111
rect 468 109 469 111
rect 465 108 469 109
rect 505 104 509 130
rect 565 132 609 133
rect 565 130 606 132
rect 608 130 609 132
rect 565 128 566 130
rect 568 129 609 130
rect 568 128 569 129
rect 565 126 569 128
rect 617 120 621 137
rect 702 138 706 139
rect 702 136 703 138
rect 705 136 706 138
rect 617 118 618 120
rect 620 118 621 120
rect 665 130 669 131
rect 665 128 666 130
rect 668 128 669 130
rect 665 122 669 128
rect 665 120 666 122
rect 668 120 669 122
rect 665 119 669 120
rect 702 119 706 136
rect 617 117 621 118
rect 702 117 703 119
rect 705 117 706 119
rect 702 116 706 117
rect 796 119 800 145
rect 796 117 797 119
rect 799 117 800 119
rect 796 116 800 117
rect 525 112 698 113
rect 525 110 526 112
rect 528 110 695 112
rect 697 110 698 112
rect 525 109 698 110
rect 804 107 808 186
rect 812 156 816 157
rect 812 154 813 156
rect 815 154 816 156
rect 812 119 816 154
rect 812 117 813 119
rect 815 117 816 119
rect 812 116 816 117
rect 725 106 808 107
rect 725 104 726 106
rect 728 104 808 106
rect 63 100 64 102
rect 66 100 67 102
rect 163 103 211 104
rect 163 101 164 103
rect 166 101 208 103
rect 210 101 211 103
rect 163 100 211 101
rect 223 103 605 104
rect 725 103 808 104
rect 223 101 224 103
rect 226 101 602 103
rect 604 101 605 103
rect 223 100 605 101
rect 63 99 67 100
rect 765 98 769 99
rect 765 96 766 98
rect 768 96 769 98
rect 24 94 730 95
rect 24 92 25 94
rect 27 92 124 94
rect 126 92 224 94
rect 226 92 324 94
rect 326 92 426 94
rect 428 92 527 94
rect 529 92 627 94
rect 629 92 727 94
rect 729 92 730 94
rect 24 91 730 92
rect 7 88 11 89
rect 7 86 8 88
rect 10 86 11 88
rect 7 37 11 86
rect 403 86 609 87
rect 403 84 404 86
rect 406 84 606 86
rect 608 84 609 86
rect 403 83 609 84
rect 765 78 769 96
rect 79 74 769 78
rect 79 54 83 74
rect 179 69 606 70
rect 179 67 466 69
rect 468 67 606 69
rect 179 66 606 67
rect 179 62 183 66
rect 602 62 606 66
rect 179 60 180 62
rect 182 60 183 62
rect 179 59 183 60
rect 279 61 506 62
rect 279 59 280 61
rect 282 59 503 61
rect 505 59 506 61
rect 602 60 603 62
rect 605 60 606 62
rect 602 59 606 60
rect 703 61 707 74
rect 703 59 704 61
rect 706 59 707 61
rect 279 58 506 59
rect 703 58 707 59
rect 79 52 80 54
rect 82 52 83 54
rect 79 51 83 52
rect 87 53 824 54
rect 87 51 88 53
rect 90 51 188 53
rect 190 51 288 53
rect 290 51 388 53
rect 390 51 488 53
rect 490 51 588 53
rect 590 51 688 53
rect 690 51 788 53
rect 790 51 821 53
rect 823 51 824 53
rect 87 50 824 51
rect 207 45 211 46
rect 207 43 208 45
rect 210 43 211 45
rect 7 35 8 37
rect 10 35 11 37
rect 7 9 11 35
rect 107 38 111 39
rect 107 36 108 38
rect 110 36 111 38
rect 107 17 111 36
rect 207 37 211 43
rect 303 45 483 46
rect 303 43 304 45
rect 306 43 308 45
rect 310 43 483 45
rect 303 42 480 43
rect 479 41 480 42
rect 482 41 483 43
rect 507 45 611 46
rect 507 43 508 45
rect 510 43 611 45
rect 507 42 611 43
rect 479 40 483 41
rect 607 38 611 42
rect 207 35 208 37
rect 210 35 211 37
rect 207 25 211 35
rect 387 37 411 38
rect 387 35 388 37
rect 390 35 404 37
rect 406 35 408 37
rect 410 35 411 37
rect 387 34 411 35
rect 587 37 591 38
rect 587 35 588 37
rect 590 35 591 37
rect 587 25 591 35
rect 607 37 669 38
rect 607 35 666 37
rect 668 35 669 37
rect 607 34 669 35
rect 687 37 691 38
rect 687 35 688 37
rect 690 35 691 37
rect 207 21 591 25
rect 687 17 691 35
rect 107 16 691 17
rect 107 14 352 16
rect 354 14 691 16
rect 107 13 691 14
rect 787 37 791 38
rect 787 35 788 37
rect 790 35 791 37
rect 787 9 791 35
rect 7 5 791 9
<< alu3 >>
rect 820 341 824 342
rect 820 339 821 341
rect 823 339 824 341
rect 200 334 443 338
rect 139 315 143 316
rect 139 313 140 315
rect 142 313 143 315
rect 30 304 34 305
rect 30 302 31 304
rect 33 302 34 304
rect 30 285 34 302
rect 30 281 104 285
rect 100 235 104 281
rect 139 252 143 313
rect 200 272 204 334
rect 299 329 304 330
rect 299 327 300 329
rect 302 327 304 329
rect 299 326 304 327
rect 200 270 201 272
rect 203 270 204 272
rect 200 269 204 270
rect 300 272 304 326
rect 439 325 443 334
rect 439 323 440 325
rect 442 323 443 325
rect 439 322 443 323
rect 598 333 602 334
rect 598 331 599 333
rect 601 331 602 333
rect 339 320 343 321
rect 339 318 340 320
rect 342 318 343 320
rect 339 288 343 318
rect 339 286 340 288
rect 342 286 343 288
rect 339 285 343 286
rect 300 270 301 272
rect 303 270 304 272
rect 300 269 304 270
rect 497 264 501 265
rect 497 262 498 264
rect 500 262 501 264
rect 497 252 501 262
rect 598 256 602 331
rect 598 254 599 256
rect 601 254 602 256
rect 598 253 602 254
rect 639 328 643 329
rect 639 326 640 328
rect 642 326 643 328
rect 139 248 501 252
rect 639 237 643 326
rect 730 304 792 305
rect 730 302 731 304
rect 733 302 792 304
rect 730 301 792 302
rect 702 288 706 289
rect 702 286 703 288
rect 705 286 706 288
rect 702 272 706 286
rect 702 270 703 272
rect 705 270 706 272
rect 702 269 706 270
rect 788 256 792 301
rect 788 254 789 256
rect 791 254 792 256
rect 788 253 792 254
rect 100 233 101 235
rect 103 233 104 235
rect 480 233 643 237
rect 100 232 104 233
rect 402 232 406 233
rect 402 230 403 232
rect 405 230 406 232
rect 402 227 406 230
rect 480 227 484 233
rect 402 223 484 227
rect 502 228 506 229
rect 502 226 503 228
rect 505 226 506 228
rect 202 222 268 223
rect 202 220 265 222
rect 267 220 268 222
rect 202 219 268 220
rect 202 181 206 219
rect 402 208 406 209
rect 402 206 403 208
rect 405 206 406 208
rect 402 189 406 206
rect 402 187 403 189
rect 405 187 406 189
rect 402 186 406 187
rect 502 189 506 226
rect 566 228 705 229
rect 566 226 567 228
rect 569 226 705 228
rect 566 225 705 226
rect 502 187 503 189
rect 505 187 506 189
rect 502 186 506 187
rect 602 220 670 221
rect 602 218 667 220
rect 669 218 670 220
rect 602 217 670 218
rect 202 179 203 181
rect 205 179 206 181
rect 202 178 206 179
rect 602 181 606 217
rect 701 189 705 225
rect 766 221 816 222
rect 766 219 767 221
rect 769 219 813 221
rect 815 219 816 221
rect 766 218 816 219
rect 701 187 702 189
rect 704 187 705 189
rect 701 186 705 187
rect 602 179 603 181
rect 605 179 606 181
rect 602 178 606 179
rect 199 166 203 167
rect 199 164 200 166
rect 202 164 203 166
rect 95 156 99 157
rect 95 154 96 156
rect 98 154 99 156
rect 95 137 99 154
rect 199 140 203 164
rect 199 138 200 140
rect 202 138 203 140
rect 199 137 203 138
rect 299 166 303 167
rect 299 164 300 166
rect 302 164 303 166
rect 95 135 96 137
rect 98 135 99 137
rect 95 134 99 135
rect 299 133 303 164
rect 402 166 501 167
rect 402 164 403 166
rect 405 164 501 166
rect 402 163 501 164
rect 497 140 501 163
rect 702 166 706 167
rect 702 164 703 166
rect 705 164 706 166
rect 497 138 498 140
rect 500 138 501 140
rect 497 137 501 138
rect 574 156 578 157
rect 574 154 575 156
rect 577 154 578 156
rect 299 132 509 133
rect 299 130 506 132
rect 508 130 509 132
rect 299 129 509 130
rect 263 123 267 124
rect 263 121 264 123
rect 266 121 267 123
rect 263 112 267 121
rect 574 120 578 154
rect 702 138 706 164
rect 774 156 816 157
rect 774 154 775 156
rect 777 154 813 156
rect 815 154 816 156
rect 774 153 816 154
rect 702 136 703 138
rect 705 136 706 138
rect 702 135 706 136
rect 295 119 578 120
rect 295 117 300 119
rect 302 117 578 119
rect 295 116 578 117
rect 605 132 609 133
rect 605 130 606 132
rect 608 130 609 132
rect 263 108 307 112
rect 207 103 211 104
rect 63 102 67 103
rect 63 100 64 102
rect 66 100 67 102
rect 63 89 67 100
rect 7 88 67 89
rect 7 86 8 88
rect 10 86 67 88
rect 7 85 67 86
rect 207 101 208 103
rect 210 101 211 103
rect 207 45 211 101
rect 207 43 208 45
rect 210 43 211 45
rect 207 42 211 43
rect 303 45 307 108
rect 303 43 304 45
rect 306 43 307 45
rect 303 42 307 43
rect 351 111 355 112
rect 351 109 352 111
rect 354 109 355 111
rect 351 16 355 109
rect 465 111 469 112
rect 465 109 466 111
rect 468 109 469 111
rect 403 86 407 87
rect 403 84 404 86
rect 406 84 407 86
rect 403 37 407 84
rect 465 69 469 109
rect 605 86 609 130
rect 605 84 606 86
rect 608 84 609 86
rect 605 83 609 84
rect 665 122 669 124
rect 665 120 666 122
rect 668 120 669 122
rect 465 67 466 69
rect 468 67 469 69
rect 465 66 469 67
rect 403 35 404 37
rect 406 35 407 37
rect 403 34 407 35
rect 665 37 669 120
rect 820 53 824 339
rect 820 51 821 53
rect 823 51 824 53
rect 820 50 824 51
rect 665 35 666 37
rect 668 35 669 37
rect 665 34 669 35
rect 351 14 352 16
rect 354 14 355 16
rect 351 13 355 14
<< ptie >>
rect 8 360 21 362
rect 8 358 10 360
rect 12 358 17 360
rect 19 358 21 360
rect 8 356 21 358
rect 108 360 121 362
rect 108 358 110 360
rect 112 358 117 360
rect 119 358 121 360
rect 108 356 121 358
rect 208 360 221 362
rect 208 358 210 360
rect 212 358 217 360
rect 219 358 221 360
rect 208 356 221 358
rect 308 360 321 362
rect 308 358 310 360
rect 312 358 317 360
rect 319 358 321 360
rect 308 356 321 358
rect 408 360 421 362
rect 408 358 410 360
rect 412 358 417 360
rect 419 358 421 360
rect 408 356 421 358
rect 508 360 521 362
rect 508 358 510 360
rect 512 358 517 360
rect 519 358 521 360
rect 508 356 521 358
rect 608 360 621 362
rect 608 358 610 360
rect 612 358 617 360
rect 619 358 621 360
rect 608 356 621 358
rect 708 360 721 362
rect 708 358 710 360
rect 712 358 717 360
rect 719 358 721 360
rect 708 356 721 358
rect 85 228 98 230
rect 85 226 87 228
rect 89 226 94 228
rect 96 226 98 228
rect 85 224 98 226
rect 185 228 198 230
rect 185 226 187 228
rect 189 226 194 228
rect 196 226 198 228
rect 185 224 198 226
rect 285 228 298 230
rect 285 226 287 228
rect 289 226 294 228
rect 296 226 298 228
rect 285 224 298 226
rect 385 228 398 230
rect 385 226 387 228
rect 389 226 394 228
rect 396 226 398 228
rect 385 224 398 226
rect 487 228 500 230
rect 487 226 489 228
rect 491 226 496 228
rect 498 226 500 228
rect 487 224 500 226
rect 587 228 600 230
rect 587 226 589 228
rect 591 226 596 228
rect 598 226 600 228
rect 587 224 600 226
rect 687 228 700 230
rect 687 226 689 228
rect 691 226 696 228
rect 698 226 700 228
rect 687 224 700 226
rect 787 228 800 230
rect 787 226 789 228
rect 791 226 796 228
rect 798 226 800 228
rect 787 224 800 226
rect 85 216 98 218
rect 85 214 87 216
rect 89 214 94 216
rect 96 214 98 216
rect 85 212 98 214
rect 185 216 198 218
rect 185 214 187 216
rect 189 214 194 216
rect 196 214 198 216
rect 185 212 198 214
rect 285 216 298 218
rect 285 214 287 216
rect 289 214 294 216
rect 296 214 298 216
rect 285 212 298 214
rect 385 216 398 218
rect 385 214 387 216
rect 389 214 394 216
rect 396 214 398 216
rect 385 212 398 214
rect 487 216 500 218
rect 487 214 489 216
rect 491 214 496 216
rect 498 214 500 216
rect 487 212 500 214
rect 587 216 600 218
rect 587 214 589 216
rect 591 214 596 216
rect 598 214 600 216
rect 587 212 600 214
rect 687 216 700 218
rect 687 214 689 216
rect 691 214 696 216
rect 698 214 700 216
rect 687 212 700 214
rect 787 216 800 218
rect 787 214 789 216
rect 791 214 796 216
rect 798 214 800 216
rect 787 212 800 214
rect 85 84 98 86
rect 85 82 87 84
rect 89 82 94 84
rect 96 82 98 84
rect 85 80 98 82
rect 185 84 198 86
rect 185 82 187 84
rect 189 82 194 84
rect 196 82 198 84
rect 185 80 198 82
rect 285 84 298 86
rect 285 82 287 84
rect 289 82 294 84
rect 296 82 298 84
rect 285 80 298 82
rect 385 84 398 86
rect 385 82 387 84
rect 389 82 394 84
rect 396 82 398 84
rect 385 80 398 82
rect 487 84 500 86
rect 487 82 489 84
rect 491 82 496 84
rect 498 82 500 84
rect 487 80 500 82
rect 587 84 600 86
rect 587 82 589 84
rect 591 82 596 84
rect 598 82 600 84
rect 587 80 600 82
rect 687 84 700 86
rect 687 82 689 84
rect 691 82 696 84
rect 698 82 700 84
rect 687 80 700 82
rect 787 84 800 86
rect 787 82 789 84
rect 791 82 796 84
rect 798 82 800 84
rect 787 80 800 82
rect 8 72 21 74
rect 8 70 10 72
rect 12 70 17 72
rect 19 70 21 72
rect 8 68 21 70
rect 108 72 121 74
rect 108 70 110 72
rect 112 70 117 72
rect 119 70 121 72
rect 108 68 121 70
rect 208 72 221 74
rect 208 70 210 72
rect 212 70 217 72
rect 219 70 221 72
rect 208 68 221 70
rect 308 72 321 74
rect 308 70 310 72
rect 312 70 317 72
rect 319 70 321 72
rect 308 68 321 70
rect 408 72 421 74
rect 408 70 410 72
rect 412 70 417 72
rect 419 70 421 72
rect 408 68 421 70
rect 508 72 521 74
rect 508 70 510 72
rect 512 70 517 72
rect 519 70 521 72
rect 508 68 521 70
rect 608 72 621 74
rect 608 70 610 72
rect 612 70 617 72
rect 619 70 621 72
rect 608 68 621 70
rect 708 72 721 74
rect 708 70 710 72
rect 712 70 717 72
rect 719 70 721 72
rect 708 68 721 70
<< ntie >>
rect 8 300 14 302
rect 8 298 10 300
rect 12 298 14 300
rect 8 296 14 298
rect 108 300 114 302
rect 108 298 110 300
rect 112 298 114 300
rect 108 296 114 298
rect 208 300 214 302
rect 208 298 210 300
rect 212 298 214 300
rect 208 296 214 298
rect 308 300 314 302
rect 308 298 310 300
rect 312 298 314 300
rect 308 296 314 298
rect 408 300 414 302
rect 408 298 410 300
rect 412 298 414 300
rect 408 296 414 298
rect 508 300 514 302
rect 508 298 510 300
rect 512 298 514 300
rect 508 296 514 298
rect 608 300 614 302
rect 608 298 610 300
rect 612 298 614 300
rect 608 296 614 298
rect 708 300 714 302
rect 708 298 710 300
rect 712 298 714 300
rect 708 296 714 298
rect 92 288 98 290
rect 92 286 94 288
rect 96 286 98 288
rect 92 284 98 286
rect 192 288 198 290
rect 192 286 194 288
rect 196 286 198 288
rect 192 284 198 286
rect 292 288 298 290
rect 292 286 294 288
rect 296 286 298 288
rect 292 284 298 286
rect 392 288 398 290
rect 392 286 394 288
rect 396 286 398 288
rect 392 284 398 286
rect 494 288 500 290
rect 494 286 496 288
rect 498 286 500 288
rect 494 284 500 286
rect 594 288 600 290
rect 594 286 596 288
rect 598 286 600 288
rect 594 284 600 286
rect 694 288 700 290
rect 694 286 696 288
rect 698 286 700 288
rect 694 284 700 286
rect 794 288 800 290
rect 794 286 796 288
rect 798 286 800 288
rect 794 284 800 286
rect 92 156 98 158
rect 92 154 94 156
rect 96 154 98 156
rect 92 152 98 154
rect 192 156 198 158
rect 192 154 194 156
rect 196 154 198 156
rect 192 152 198 154
rect 292 156 298 158
rect 292 154 294 156
rect 296 154 298 156
rect 292 152 298 154
rect 392 156 398 158
rect 392 154 394 156
rect 396 154 398 156
rect 392 152 398 154
rect 494 156 500 158
rect 494 154 496 156
rect 498 154 500 156
rect 494 152 500 154
rect 594 156 600 158
rect 594 154 596 156
rect 598 154 600 156
rect 594 152 600 154
rect 694 156 700 158
rect 694 154 696 156
rect 698 154 700 156
rect 694 152 700 154
rect 794 156 800 158
rect 794 154 796 156
rect 798 154 800 156
rect 794 152 800 154
rect 92 144 98 146
rect 92 142 94 144
rect 96 142 98 144
rect 92 140 98 142
rect 192 144 198 146
rect 192 142 194 144
rect 196 142 198 144
rect 192 140 198 142
rect 292 144 298 146
rect 292 142 294 144
rect 296 142 298 144
rect 292 140 298 142
rect 392 144 398 146
rect 392 142 394 144
rect 396 142 398 144
rect 392 140 398 142
rect 494 144 500 146
rect 494 142 496 144
rect 498 142 500 144
rect 494 140 500 142
rect 594 144 600 146
rect 594 142 596 144
rect 598 142 600 144
rect 594 140 600 142
rect 694 144 700 146
rect 694 142 696 144
rect 698 142 700 144
rect 694 140 700 142
rect 794 144 800 146
rect 794 142 796 144
rect 798 142 800 144
rect 794 140 800 142
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 108 12 114 14
rect 108 10 110 12
rect 112 10 114 12
rect 108 8 114 10
rect 208 12 214 14
rect 208 10 210 12
rect 212 10 214 12
rect 208 8 214 10
rect 308 12 314 14
rect 308 10 310 12
rect 312 10 314 12
rect 308 8 314 10
rect 408 12 414 14
rect 408 10 410 12
rect 412 10 414 12
rect 408 8 414 10
rect 508 12 514 14
rect 508 10 510 12
rect 512 10 514 12
rect 508 8 514 10
rect 608 12 614 14
rect 608 10 610 12
rect 612 10 614 12
rect 608 8 614 10
rect 708 12 714 14
rect 708 10 710 12
rect 712 10 714 12
rect 708 8 714 10
<< nmos >>
rect 16 340 18 350
rect 27 340 29 351
rect 37 340 39 351
rect 47 345 49 356
rect 57 342 59 353
rect 77 342 79 352
rect 90 342 92 349
rect 116 340 118 350
rect 127 340 129 351
rect 137 340 139 351
rect 147 345 149 356
rect 157 342 159 353
rect 177 342 179 352
rect 190 342 192 349
rect 216 340 218 350
rect 227 340 229 351
rect 237 340 239 351
rect 247 345 249 356
rect 257 342 259 353
rect 277 342 279 352
rect 290 342 292 349
rect 316 340 318 350
rect 327 340 329 351
rect 337 340 339 351
rect 347 345 349 356
rect 357 342 359 353
rect 377 342 379 352
rect 390 342 392 349
rect 416 340 418 350
rect 427 340 429 351
rect 437 340 439 351
rect 447 345 449 356
rect 457 342 459 353
rect 477 342 479 352
rect 490 342 492 349
rect 516 340 518 350
rect 527 340 529 351
rect 537 340 539 351
rect 547 345 549 356
rect 557 342 559 353
rect 577 342 579 352
rect 590 342 592 349
rect 616 340 618 350
rect 627 340 629 351
rect 637 340 639 351
rect 647 345 649 356
rect 657 342 659 353
rect 677 342 679 352
rect 690 342 692 349
rect 716 340 718 350
rect 727 340 729 351
rect 737 340 739 351
rect 747 345 749 356
rect 757 342 759 353
rect 777 342 779 352
rect 790 342 792 349
rect 14 237 16 244
rect 27 234 29 244
rect 47 233 49 244
rect 57 230 59 241
rect 67 235 69 246
rect 77 235 79 246
rect 88 236 90 246
rect 114 237 116 244
rect 127 234 129 244
rect 147 233 149 244
rect 157 230 159 241
rect 167 235 169 246
rect 177 235 179 246
rect 188 236 190 246
rect 214 237 216 244
rect 227 234 229 244
rect 247 233 249 244
rect 257 230 259 241
rect 267 235 269 246
rect 277 235 279 246
rect 288 236 290 246
rect 314 237 316 244
rect 327 234 329 244
rect 347 233 349 244
rect 357 230 359 241
rect 367 235 369 246
rect 377 235 379 246
rect 388 236 390 246
rect 416 237 418 244
rect 429 234 431 244
rect 449 233 451 244
rect 459 230 461 241
rect 469 235 471 246
rect 479 235 481 246
rect 490 236 492 246
rect 516 237 518 244
rect 529 234 531 244
rect 549 233 551 244
rect 559 230 561 241
rect 569 235 571 246
rect 579 235 581 246
rect 590 236 592 246
rect 616 237 618 244
rect 629 234 631 244
rect 649 233 651 244
rect 659 230 661 241
rect 669 235 671 246
rect 679 235 681 246
rect 690 236 692 246
rect 716 237 718 244
rect 729 234 731 244
rect 749 233 751 244
rect 759 230 761 241
rect 769 235 771 246
rect 779 235 781 246
rect 790 236 792 246
rect 14 198 16 205
rect 27 198 29 208
rect 47 198 49 209
rect 57 201 59 212
rect 67 196 69 207
rect 77 196 79 207
rect 88 196 90 206
rect 114 198 116 205
rect 127 198 129 208
rect 147 198 149 209
rect 157 201 159 212
rect 167 196 169 207
rect 177 196 179 207
rect 188 196 190 206
rect 214 198 216 205
rect 227 198 229 208
rect 247 198 249 209
rect 257 201 259 212
rect 267 196 269 207
rect 277 196 279 207
rect 288 196 290 206
rect 314 198 316 205
rect 327 198 329 208
rect 347 198 349 209
rect 357 201 359 212
rect 367 196 369 207
rect 377 196 379 207
rect 388 196 390 206
rect 416 198 418 205
rect 429 198 431 208
rect 449 198 451 209
rect 459 201 461 212
rect 469 196 471 207
rect 479 196 481 207
rect 490 196 492 206
rect 516 198 518 205
rect 529 198 531 208
rect 549 198 551 209
rect 559 201 561 212
rect 569 196 571 207
rect 579 196 581 207
rect 590 196 592 206
rect 616 198 618 205
rect 629 198 631 208
rect 649 198 651 209
rect 659 201 661 212
rect 669 196 671 207
rect 679 196 681 207
rect 690 196 692 206
rect 716 198 718 205
rect 729 198 731 208
rect 749 198 751 209
rect 759 201 761 212
rect 769 196 771 207
rect 779 196 781 207
rect 790 196 792 206
rect 14 93 16 100
rect 27 90 29 100
rect 47 89 49 100
rect 57 86 59 97
rect 67 91 69 102
rect 77 91 79 102
rect 88 92 90 102
rect 114 93 116 100
rect 127 90 129 100
rect 147 89 149 100
rect 157 86 159 97
rect 167 91 169 102
rect 177 91 179 102
rect 188 92 190 102
rect 214 93 216 100
rect 227 90 229 100
rect 247 89 249 100
rect 257 86 259 97
rect 267 91 269 102
rect 277 91 279 102
rect 288 92 290 102
rect 314 93 316 100
rect 327 90 329 100
rect 347 89 349 100
rect 357 86 359 97
rect 367 91 369 102
rect 377 91 379 102
rect 388 92 390 102
rect 416 93 418 100
rect 429 90 431 100
rect 449 89 451 100
rect 459 86 461 97
rect 469 91 471 102
rect 479 91 481 102
rect 490 92 492 102
rect 516 93 518 100
rect 529 90 531 100
rect 549 89 551 100
rect 559 86 561 97
rect 569 91 571 102
rect 579 91 581 102
rect 590 92 592 102
rect 616 93 618 100
rect 629 90 631 100
rect 649 89 651 100
rect 659 86 661 97
rect 669 91 671 102
rect 679 91 681 102
rect 690 92 692 102
rect 716 93 718 100
rect 729 90 731 100
rect 749 89 751 100
rect 759 86 761 97
rect 769 91 771 102
rect 779 91 781 102
rect 790 92 792 102
rect 16 52 18 62
rect 27 52 29 63
rect 37 52 39 63
rect 47 57 49 68
rect 57 54 59 65
rect 77 54 79 64
rect 90 54 92 61
rect 116 52 118 62
rect 127 52 129 63
rect 137 52 139 63
rect 147 57 149 68
rect 157 54 159 65
rect 177 54 179 64
rect 190 54 192 61
rect 216 52 218 62
rect 227 52 229 63
rect 237 52 239 63
rect 247 57 249 68
rect 257 54 259 65
rect 277 54 279 64
rect 290 54 292 61
rect 316 52 318 62
rect 327 52 329 63
rect 337 52 339 63
rect 347 57 349 68
rect 357 54 359 65
rect 377 54 379 64
rect 390 54 392 61
rect 416 52 418 62
rect 427 52 429 63
rect 437 52 439 63
rect 447 57 449 68
rect 457 54 459 65
rect 477 54 479 64
rect 490 54 492 61
rect 516 52 518 62
rect 527 52 529 63
rect 537 52 539 63
rect 547 57 549 68
rect 557 54 559 65
rect 577 54 579 64
rect 590 54 592 61
rect 616 52 618 62
rect 627 52 629 63
rect 637 52 639 63
rect 647 57 649 68
rect 657 54 659 65
rect 677 54 679 64
rect 690 54 692 61
rect 716 52 718 62
rect 727 52 729 63
rect 737 52 739 63
rect 747 57 749 68
rect 757 54 759 65
rect 777 54 779 64
rect 790 54 792 61
<< pmos >>
rect 14 314 16 327
rect 25 305 27 327
rect 35 305 37 327
rect 45 305 47 327
rect 59 305 61 327
rect 77 314 79 327
rect 90 309 92 319
rect 114 314 116 327
rect 125 305 127 327
rect 135 305 137 327
rect 145 305 147 327
rect 159 305 161 327
rect 177 314 179 327
rect 190 309 192 319
rect 214 314 216 327
rect 225 305 227 327
rect 235 305 237 327
rect 245 305 247 327
rect 259 305 261 327
rect 277 314 279 327
rect 290 309 292 319
rect 314 314 316 327
rect 325 305 327 327
rect 335 305 337 327
rect 345 305 347 327
rect 359 305 361 327
rect 377 314 379 327
rect 390 309 392 319
rect 414 314 416 327
rect 425 305 427 327
rect 435 305 437 327
rect 445 305 447 327
rect 459 305 461 327
rect 477 314 479 327
rect 490 309 492 319
rect 514 314 516 327
rect 525 305 527 327
rect 535 305 537 327
rect 545 305 547 327
rect 559 305 561 327
rect 577 314 579 327
rect 590 309 592 319
rect 614 314 616 327
rect 625 305 627 327
rect 635 305 637 327
rect 645 305 647 327
rect 659 305 661 327
rect 677 314 679 327
rect 690 309 692 319
rect 714 314 716 327
rect 725 305 727 327
rect 735 305 737 327
rect 745 305 747 327
rect 759 305 761 327
rect 777 314 779 327
rect 790 309 792 319
rect 14 267 16 277
rect 27 259 29 272
rect 45 259 47 281
rect 59 259 61 281
rect 69 259 71 281
rect 79 259 81 281
rect 90 259 92 272
rect 114 267 116 277
rect 127 259 129 272
rect 145 259 147 281
rect 159 259 161 281
rect 169 259 171 281
rect 179 259 181 281
rect 190 259 192 272
rect 214 267 216 277
rect 227 259 229 272
rect 245 259 247 281
rect 259 259 261 281
rect 269 259 271 281
rect 279 259 281 281
rect 290 259 292 273
rect 314 267 316 277
rect 327 259 329 272
rect 345 259 347 281
rect 359 259 361 281
rect 369 259 371 281
rect 379 259 381 281
rect 390 259 392 272
rect 416 267 418 277
rect 429 259 431 272
rect 447 259 449 281
rect 461 259 463 281
rect 471 259 473 281
rect 481 259 483 281
rect 492 260 494 273
rect 516 267 518 277
rect 529 259 531 272
rect 547 259 549 281
rect 561 259 563 281
rect 571 259 573 281
rect 581 259 583 281
rect 592 259 594 272
rect 616 267 618 277
rect 629 259 631 272
rect 647 259 649 281
rect 661 259 663 281
rect 671 259 673 281
rect 681 259 683 281
rect 692 260 694 273
rect 716 267 718 277
rect 729 259 731 272
rect 747 259 749 281
rect 761 259 763 281
rect 771 259 773 281
rect 781 259 783 281
rect 792 259 794 272
rect 14 165 16 175
rect 27 170 29 183
rect 45 161 47 183
rect 59 161 61 183
rect 69 161 71 183
rect 79 161 81 183
rect 90 170 92 183
rect 114 165 116 175
rect 127 170 129 183
rect 145 161 147 183
rect 159 161 161 183
rect 169 161 171 183
rect 179 161 181 183
rect 190 170 192 183
rect 214 165 216 175
rect 227 170 229 183
rect 245 161 247 183
rect 259 161 261 183
rect 269 161 271 183
rect 279 161 281 183
rect 290 170 292 183
rect 314 165 316 175
rect 327 170 329 183
rect 345 161 347 183
rect 359 161 361 183
rect 369 161 371 183
rect 379 161 381 183
rect 390 170 392 183
rect 416 165 418 175
rect 429 170 431 183
rect 447 161 449 183
rect 461 161 463 183
rect 471 161 473 183
rect 481 161 483 183
rect 492 170 494 183
rect 516 165 518 175
rect 529 170 531 183
rect 547 161 549 183
rect 561 161 563 183
rect 571 161 573 183
rect 581 161 583 183
rect 592 170 594 183
rect 616 165 618 175
rect 629 170 631 183
rect 647 161 649 183
rect 661 161 663 183
rect 671 161 673 183
rect 681 161 683 183
rect 692 170 694 183
rect 716 165 718 175
rect 729 170 731 183
rect 747 161 749 183
rect 761 161 763 183
rect 771 161 773 183
rect 781 161 783 183
rect 792 170 794 183
rect 14 123 16 133
rect 27 115 29 128
rect 45 115 47 137
rect 59 115 61 137
rect 69 115 71 137
rect 79 115 81 137
rect 90 115 92 128
rect 114 123 116 133
rect 127 115 129 128
rect 145 115 147 137
rect 159 115 161 137
rect 169 115 171 137
rect 179 115 181 137
rect 190 115 192 128
rect 214 123 216 133
rect 227 115 229 128
rect 245 115 247 137
rect 259 115 261 137
rect 269 115 271 137
rect 279 115 281 137
rect 290 115 292 128
rect 314 123 316 133
rect 327 115 329 128
rect 345 115 347 137
rect 359 115 361 137
rect 369 115 371 137
rect 379 115 381 137
rect 390 115 392 128
rect 416 123 418 133
rect 429 115 431 128
rect 447 115 449 137
rect 461 115 463 137
rect 471 115 473 137
rect 481 115 483 137
rect 492 115 494 128
rect 516 123 518 133
rect 529 115 531 128
rect 547 115 549 137
rect 561 115 563 137
rect 571 115 573 137
rect 581 115 583 137
rect 592 115 594 128
rect 616 123 618 133
rect 629 115 631 128
rect 647 115 649 137
rect 661 115 663 137
rect 671 115 673 137
rect 681 115 683 137
rect 692 115 694 128
rect 716 123 718 133
rect 729 115 731 128
rect 747 115 749 137
rect 761 115 763 137
rect 771 115 773 137
rect 781 115 783 137
rect 792 115 794 128
rect 14 26 16 39
rect 25 17 27 39
rect 35 17 37 39
rect 45 17 47 39
rect 59 17 61 39
rect 77 26 79 39
rect 90 21 92 31
rect 114 26 116 39
rect 125 17 127 39
rect 135 17 137 39
rect 145 17 147 39
rect 159 17 161 39
rect 177 26 179 39
rect 190 21 192 31
rect 214 26 216 39
rect 225 17 227 39
rect 235 17 237 39
rect 245 17 247 39
rect 259 17 261 39
rect 277 26 279 39
rect 290 21 292 31
rect 314 26 316 39
rect 325 17 327 39
rect 335 17 337 39
rect 345 17 347 39
rect 359 17 361 39
rect 377 26 379 39
rect 390 21 392 31
rect 414 26 416 39
rect 425 17 427 39
rect 435 17 437 39
rect 445 17 447 39
rect 459 17 461 39
rect 477 26 479 39
rect 490 21 492 31
rect 514 26 516 39
rect 525 17 527 39
rect 535 17 537 39
rect 545 17 547 39
rect 559 17 561 39
rect 577 26 579 39
rect 590 21 592 31
rect 614 26 616 39
rect 625 17 627 39
rect 635 17 637 39
rect 645 17 647 39
rect 659 17 661 39
rect 677 26 679 39
rect 690 21 692 31
rect 714 26 716 39
rect 725 17 727 39
rect 735 17 737 39
rect 745 17 747 39
rect 759 17 761 39
rect 777 26 779 39
rect 790 21 792 31
<< polyct0 >>
rect 25 332 27 334
rect 47 332 49 334
rect 62 332 64 334
rect 125 332 127 334
rect 147 332 149 334
rect 162 332 164 334
rect 225 332 227 334
rect 247 332 249 334
rect 262 332 264 334
rect 325 332 327 334
rect 347 332 349 334
rect 362 332 364 334
rect 425 332 427 334
rect 447 332 449 334
rect 462 332 464 334
rect 525 332 527 334
rect 547 332 549 334
rect 562 332 564 334
rect 625 332 627 334
rect 647 332 649 334
rect 662 332 664 334
rect 725 332 727 334
rect 747 332 749 334
rect 762 332 764 334
rect 42 252 44 254
rect 57 252 59 254
rect 79 252 81 254
rect 142 252 144 254
rect 157 252 159 254
rect 179 252 181 254
rect 242 252 244 254
rect 257 252 259 254
rect 279 252 281 254
rect 342 252 344 254
rect 357 252 359 254
rect 379 252 381 254
rect 444 252 446 254
rect 459 252 461 254
rect 481 252 483 254
rect 544 252 546 254
rect 559 252 561 254
rect 581 252 583 254
rect 644 252 646 254
rect 659 252 661 254
rect 681 252 683 254
rect 744 252 746 254
rect 759 252 761 254
rect 781 252 783 254
rect 42 188 44 190
rect 57 188 59 190
rect 79 188 81 190
rect 142 188 144 190
rect 157 188 159 190
rect 179 188 181 190
rect 242 188 244 190
rect 257 188 259 190
rect 279 188 281 190
rect 342 188 344 190
rect 357 188 359 190
rect 379 188 381 190
rect 444 188 446 190
rect 459 188 461 190
rect 481 188 483 190
rect 544 188 546 190
rect 559 188 561 190
rect 581 188 583 190
rect 644 188 646 190
rect 659 188 661 190
rect 681 188 683 190
rect 744 188 746 190
rect 759 188 761 190
rect 781 188 783 190
rect 42 108 44 110
rect 57 108 59 110
rect 79 108 81 110
rect 142 108 144 110
rect 157 108 159 110
rect 179 108 181 110
rect 242 108 244 110
rect 257 108 259 110
rect 279 108 281 110
rect 342 108 344 110
rect 357 108 359 110
rect 379 108 381 110
rect 444 108 446 110
rect 459 108 461 110
rect 481 108 483 110
rect 544 108 546 110
rect 559 108 561 110
rect 581 108 583 110
rect 644 108 646 110
rect 659 108 661 110
rect 681 108 683 110
rect 744 108 746 110
rect 759 108 761 110
rect 781 108 783 110
rect 25 44 27 46
rect 47 44 49 46
rect 62 44 64 46
rect 125 44 127 46
rect 147 44 149 46
rect 162 44 164 46
rect 225 44 227 46
rect 247 44 249 46
rect 262 44 264 46
rect 325 44 327 46
rect 347 44 349 46
rect 362 44 364 46
rect 425 44 427 46
rect 447 44 449 46
rect 462 44 464 46
rect 525 44 527 46
rect 547 44 549 46
rect 562 44 564 46
rect 625 44 627 46
rect 647 44 649 46
rect 662 44 664 46
rect 725 44 727 46
rect 747 44 749 46
rect 762 44 764 46
<< polyct1 >>
rect 14 332 16 334
rect 78 333 80 335
rect 88 335 90 337
rect 114 332 116 334
rect 178 333 180 335
rect 188 335 190 337
rect 214 332 216 334
rect 278 333 280 335
rect 288 335 290 337
rect 314 332 316 334
rect 378 333 380 335
rect 388 335 390 337
rect 414 332 416 334
rect 478 333 480 335
rect 488 335 490 337
rect 514 332 516 334
rect 578 333 580 335
rect 588 335 590 337
rect 614 332 616 334
rect 678 333 680 335
rect 688 335 690 337
rect 714 332 716 334
rect 778 333 780 335
rect 788 335 790 337
rect 16 249 18 251
rect 26 251 28 253
rect 90 252 92 254
rect 116 249 118 251
rect 126 251 128 253
rect 190 252 192 254
rect 216 249 218 251
rect 226 251 228 253
rect 290 252 292 254
rect 316 249 318 251
rect 326 251 328 253
rect 390 252 392 254
rect 418 249 420 251
rect 428 251 430 253
rect 492 252 494 254
rect 518 249 520 251
rect 528 251 530 253
rect 592 252 594 254
rect 618 249 620 251
rect 628 251 630 253
rect 692 252 694 254
rect 718 249 720 251
rect 728 251 730 253
rect 792 252 794 254
rect 16 191 18 193
rect 26 189 28 191
rect 90 188 92 190
rect 116 191 118 193
rect 126 190 128 192
rect 190 188 192 190
rect 216 191 218 193
rect 226 189 228 191
rect 290 188 292 190
rect 316 191 318 193
rect 326 190 328 192
rect 389 188 391 190
rect 418 191 420 193
rect 428 189 430 191
rect 492 188 494 190
rect 518 191 520 193
rect 528 190 530 192
rect 592 188 594 190
rect 618 191 620 193
rect 628 189 630 191
rect 692 188 694 190
rect 718 191 720 193
rect 728 190 730 192
rect 792 188 794 190
rect 16 105 18 107
rect 26 107 28 109
rect 90 108 92 110
rect 116 105 118 107
rect 127 107 129 109
rect 190 108 192 110
rect 216 105 218 107
rect 226 107 228 109
rect 290 108 292 110
rect 316 105 318 107
rect 326 107 328 109
rect 390 108 392 110
rect 418 105 420 107
rect 428 107 430 109
rect 492 108 494 110
rect 518 105 520 107
rect 528 107 530 109
rect 592 108 594 110
rect 618 105 620 107
rect 628 107 630 109
rect 692 108 694 110
rect 718 105 720 107
rect 728 107 730 109
rect 792 108 794 110
rect 14 44 16 46
rect 78 45 80 47
rect 88 47 90 49
rect 114 44 116 46
rect 178 45 180 47
rect 188 47 190 49
rect 214 44 216 46
rect 278 45 280 47
rect 288 47 290 49
rect 314 44 316 46
rect 378 45 380 47
rect 388 47 390 49
rect 414 44 416 46
rect 478 45 480 47
rect 488 47 490 49
rect 514 44 516 46
rect 578 45 580 47
rect 588 47 590 49
rect 614 44 616 46
rect 678 45 680 47
rect 688 47 690 49
rect 714 44 716 46
rect 778 45 780 47
rect 788 47 790 49
<< ndifct0 >>
rect 11 342 13 344
rect 22 347 24 349
rect 32 342 34 344
rect 52 347 54 349
rect 84 355 86 357
rect 62 349 64 351
rect 72 344 74 346
rect 95 344 97 346
rect 111 342 113 344
rect 122 347 124 349
rect 132 342 134 344
rect 152 347 154 349
rect 184 355 186 357
rect 162 349 164 351
rect 172 344 174 346
rect 195 344 197 346
rect 211 342 213 344
rect 222 347 224 349
rect 232 342 234 344
rect 252 347 254 349
rect 284 355 286 357
rect 262 349 264 351
rect 272 344 274 346
rect 295 344 297 346
rect 311 342 313 344
rect 322 347 324 349
rect 332 342 334 344
rect 352 347 354 349
rect 384 355 386 357
rect 362 349 364 351
rect 372 344 374 346
rect 395 344 397 346
rect 411 342 413 344
rect 422 347 424 349
rect 432 342 434 344
rect 452 347 454 349
rect 484 355 486 357
rect 462 349 464 351
rect 472 344 474 346
rect 495 344 497 346
rect 511 342 513 344
rect 522 347 524 349
rect 532 342 534 344
rect 552 347 554 349
rect 584 355 586 357
rect 562 349 564 351
rect 572 344 574 346
rect 595 344 597 346
rect 611 342 613 344
rect 622 347 624 349
rect 632 342 634 344
rect 652 347 654 349
rect 684 355 686 357
rect 662 349 664 351
rect 672 344 674 346
rect 695 344 697 346
rect 711 342 713 344
rect 722 347 724 349
rect 732 342 734 344
rect 752 347 754 349
rect 784 355 786 357
rect 762 349 764 351
rect 772 344 774 346
rect 795 344 797 346
rect 9 240 11 242
rect 32 240 34 242
rect 42 235 44 237
rect 20 229 22 231
rect 52 237 54 239
rect 72 242 74 244
rect 82 237 84 239
rect 93 242 95 244
rect 109 240 111 242
rect 132 240 134 242
rect 142 235 144 237
rect 120 229 122 231
rect 152 237 154 239
rect 172 242 174 244
rect 182 237 184 239
rect 193 242 195 244
rect 209 240 211 242
rect 232 240 234 242
rect 242 235 244 237
rect 220 229 222 231
rect 252 237 254 239
rect 272 242 274 244
rect 282 237 284 239
rect 293 242 295 244
rect 309 240 311 242
rect 332 240 334 242
rect 342 235 344 237
rect 320 229 322 231
rect 352 237 354 239
rect 372 242 374 244
rect 382 237 384 239
rect 393 242 395 244
rect 411 240 413 242
rect 434 240 436 242
rect 444 235 446 237
rect 422 229 424 231
rect 454 237 456 239
rect 474 242 476 244
rect 484 237 486 239
rect 495 242 497 244
rect 511 240 513 242
rect 534 240 536 242
rect 544 235 546 237
rect 522 229 524 231
rect 554 237 556 239
rect 574 242 576 244
rect 584 237 586 239
rect 595 242 597 244
rect 611 240 613 242
rect 634 240 636 242
rect 644 235 646 237
rect 622 229 624 231
rect 654 237 656 239
rect 674 242 676 244
rect 684 237 686 239
rect 695 242 697 244
rect 711 240 713 242
rect 734 240 736 242
rect 744 235 746 237
rect 722 229 724 231
rect 754 237 756 239
rect 774 242 776 244
rect 784 237 786 239
rect 795 242 797 244
rect 20 211 22 213
rect 9 200 11 202
rect 42 205 44 207
rect 32 200 34 202
rect 52 203 54 205
rect 72 198 74 200
rect 82 203 84 205
rect 120 211 122 213
rect 93 198 95 200
rect 109 200 111 202
rect 142 205 144 207
rect 132 200 134 202
rect 152 203 154 205
rect 172 198 174 200
rect 182 203 184 205
rect 220 211 222 213
rect 193 198 195 200
rect 209 200 211 202
rect 242 205 244 207
rect 232 200 234 202
rect 252 203 254 205
rect 272 198 274 200
rect 282 203 284 205
rect 320 211 322 213
rect 293 198 295 200
rect 309 200 311 202
rect 342 205 344 207
rect 332 200 334 202
rect 352 203 354 205
rect 372 198 374 200
rect 382 203 384 205
rect 422 211 424 213
rect 393 198 395 200
rect 411 200 413 202
rect 444 205 446 207
rect 434 200 436 202
rect 454 203 456 205
rect 474 198 476 200
rect 484 203 486 205
rect 522 211 524 213
rect 495 198 497 200
rect 511 200 513 202
rect 544 205 546 207
rect 534 200 536 202
rect 554 203 556 205
rect 574 198 576 200
rect 584 203 586 205
rect 622 211 624 213
rect 595 198 597 200
rect 611 200 613 202
rect 644 205 646 207
rect 634 200 636 202
rect 654 203 656 205
rect 674 198 676 200
rect 684 203 686 205
rect 722 211 724 213
rect 695 198 697 200
rect 711 200 713 202
rect 744 205 746 207
rect 734 200 736 202
rect 754 203 756 205
rect 774 198 776 200
rect 784 203 786 205
rect 795 198 797 200
rect 9 96 11 98
rect 32 96 34 98
rect 42 91 44 93
rect 20 85 22 87
rect 52 93 54 95
rect 72 98 74 100
rect 82 93 84 95
rect 93 98 95 100
rect 109 96 111 98
rect 132 96 134 98
rect 142 91 144 93
rect 120 85 122 87
rect 152 93 154 95
rect 172 98 174 100
rect 182 93 184 95
rect 193 98 195 100
rect 209 96 211 98
rect 232 96 234 98
rect 242 91 244 93
rect 220 85 222 87
rect 252 93 254 95
rect 272 98 274 100
rect 282 93 284 95
rect 293 98 295 100
rect 309 96 311 98
rect 332 96 334 98
rect 342 91 344 93
rect 320 85 322 87
rect 352 93 354 95
rect 372 98 374 100
rect 382 93 384 95
rect 393 98 395 100
rect 411 96 413 98
rect 434 96 436 98
rect 444 91 446 93
rect 422 85 424 87
rect 454 93 456 95
rect 474 98 476 100
rect 484 93 486 95
rect 495 98 497 100
rect 511 96 513 98
rect 534 96 536 98
rect 544 91 546 93
rect 522 85 524 87
rect 554 93 556 95
rect 574 98 576 100
rect 584 93 586 95
rect 595 98 597 100
rect 611 96 613 98
rect 634 96 636 98
rect 644 91 646 93
rect 622 85 624 87
rect 654 93 656 95
rect 674 98 676 100
rect 684 93 686 95
rect 695 98 697 100
rect 711 96 713 98
rect 734 96 736 98
rect 744 91 746 93
rect 722 85 724 87
rect 754 93 756 95
rect 774 98 776 100
rect 784 93 786 95
rect 795 98 797 100
rect 11 54 13 56
rect 22 59 24 61
rect 32 54 34 56
rect 52 59 54 61
rect 84 67 86 69
rect 62 61 64 63
rect 72 56 74 58
rect 95 56 97 58
rect 111 54 113 56
rect 122 59 124 61
rect 132 54 134 56
rect 152 59 154 61
rect 184 67 186 69
rect 162 61 164 63
rect 172 56 174 58
rect 195 56 197 58
rect 211 54 213 56
rect 222 59 224 61
rect 232 54 234 56
rect 252 59 254 61
rect 284 67 286 69
rect 262 61 264 63
rect 272 56 274 58
rect 295 56 297 58
rect 311 54 313 56
rect 322 59 324 61
rect 332 54 334 56
rect 352 59 354 61
rect 384 67 386 69
rect 362 61 364 63
rect 372 56 374 58
rect 395 56 397 58
rect 411 54 413 56
rect 422 59 424 61
rect 432 54 434 56
rect 452 59 454 61
rect 484 67 486 69
rect 462 61 464 63
rect 472 56 474 58
rect 495 56 497 58
rect 511 54 513 56
rect 522 59 524 61
rect 532 54 534 56
rect 552 59 554 61
rect 584 67 586 69
rect 562 61 564 63
rect 572 56 574 58
rect 595 56 597 58
rect 611 54 613 56
rect 622 59 624 61
rect 632 54 634 56
rect 652 59 654 61
rect 684 67 686 69
rect 662 61 664 63
rect 672 56 674 58
rect 695 56 697 58
rect 711 54 713 56
rect 722 59 724 61
rect 732 54 734 56
rect 752 59 754 61
rect 784 67 786 69
rect 762 61 764 63
rect 772 56 774 58
rect 795 56 797 58
<< ndifct1 >>
rect 42 347 44 349
rect 142 347 144 349
rect 242 347 244 349
rect 342 347 344 349
rect 442 347 444 349
rect 542 347 544 349
rect 642 347 644 349
rect 742 347 744 349
rect 62 237 64 239
rect 162 237 164 239
rect 262 237 264 239
rect 362 237 364 239
rect 464 237 466 239
rect 564 237 566 239
rect 664 237 666 239
rect 764 237 766 239
rect 62 203 64 205
rect 162 203 164 205
rect 262 203 264 205
rect 362 203 364 205
rect 464 203 466 205
rect 564 203 566 205
rect 664 203 666 205
rect 764 203 766 205
rect 62 93 64 95
rect 162 93 164 95
rect 262 93 264 95
rect 362 93 364 95
rect 464 93 466 95
rect 564 93 566 95
rect 664 93 666 95
rect 764 93 766 95
rect 42 59 44 61
rect 142 59 144 61
rect 242 59 244 61
rect 342 59 344 61
rect 442 59 444 61
rect 542 59 544 61
rect 642 59 644 61
rect 742 59 744 61
<< ntiect1 >>
rect 10 298 12 300
rect 110 298 112 300
rect 210 298 212 300
rect 310 298 312 300
rect 410 298 412 300
rect 510 298 512 300
rect 610 298 612 300
rect 710 298 712 300
rect 94 286 96 288
rect 194 286 196 288
rect 294 286 296 288
rect 394 286 396 288
rect 496 286 498 288
rect 596 286 598 288
rect 696 286 698 288
rect 796 286 798 288
rect 94 154 96 156
rect 194 154 196 156
rect 294 154 296 156
rect 394 154 396 156
rect 496 154 498 156
rect 596 154 598 156
rect 696 154 698 156
rect 796 154 798 156
rect 94 142 96 144
rect 194 142 196 144
rect 294 142 296 144
rect 394 142 396 144
rect 496 142 498 144
rect 596 142 598 144
rect 696 142 698 144
rect 796 142 798 144
rect 10 10 12 12
rect 110 10 112 12
rect 210 10 212 12
rect 310 10 312 12
rect 410 10 412 12
rect 510 10 512 12
rect 610 10 612 12
rect 710 10 712 12
<< ptiect1 >>
rect 10 358 12 360
rect 17 358 19 360
rect 110 358 112 360
rect 117 358 119 360
rect 210 358 212 360
rect 217 358 219 360
rect 310 358 312 360
rect 317 358 319 360
rect 410 358 412 360
rect 417 358 419 360
rect 510 358 512 360
rect 517 358 519 360
rect 610 358 612 360
rect 617 358 619 360
rect 710 358 712 360
rect 717 358 719 360
rect 87 226 89 228
rect 94 226 96 228
rect 187 226 189 228
rect 194 226 196 228
rect 287 226 289 228
rect 294 226 296 228
rect 387 226 389 228
rect 394 226 396 228
rect 489 226 491 228
rect 496 226 498 228
rect 589 226 591 228
rect 596 226 598 228
rect 689 226 691 228
rect 696 226 698 228
rect 789 226 791 228
rect 796 226 798 228
rect 87 214 89 216
rect 94 214 96 216
rect 187 214 189 216
rect 194 214 196 216
rect 287 214 289 216
rect 294 214 296 216
rect 387 214 389 216
rect 394 214 396 216
rect 489 214 491 216
rect 496 214 498 216
rect 589 214 591 216
rect 596 214 598 216
rect 689 214 691 216
rect 696 214 698 216
rect 789 214 791 216
rect 796 214 798 216
rect 87 82 89 84
rect 94 82 96 84
rect 187 82 189 84
rect 194 82 196 84
rect 287 82 289 84
rect 294 82 296 84
rect 387 82 389 84
rect 394 82 396 84
rect 489 82 491 84
rect 496 82 498 84
rect 589 82 591 84
rect 596 82 598 84
rect 689 82 691 84
rect 696 82 698 84
rect 789 82 791 84
rect 796 82 798 84
rect 10 70 12 72
rect 17 70 19 72
rect 110 70 112 72
rect 117 70 119 72
rect 210 70 212 72
rect 217 70 219 72
rect 310 70 312 72
rect 317 70 319 72
rect 410 70 412 72
rect 417 70 419 72
rect 510 70 512 72
rect 517 70 519 72
rect 610 70 612 72
rect 617 70 619 72
rect 710 70 712 72
rect 717 70 719 72
<< pdifct0 >>
rect 9 316 11 318
rect 20 308 22 310
rect 30 316 32 318
rect 54 323 56 325
rect 72 323 74 325
rect 95 315 97 317
rect 64 307 66 309
rect 83 307 85 309
rect 120 308 122 310
rect 130 316 132 318
rect 154 323 156 325
rect 172 323 174 325
rect 195 315 197 317
rect 209 316 211 318
rect 164 307 166 309
rect 183 307 185 309
rect 220 308 222 310
rect 230 316 232 318
rect 254 323 256 325
rect 272 323 274 325
rect 295 315 297 317
rect 309 316 311 318
rect 264 307 266 309
rect 283 307 285 309
rect 320 308 322 310
rect 330 316 332 318
rect 354 323 356 325
rect 372 323 374 325
rect 395 315 397 317
rect 409 316 411 318
rect 364 307 366 309
rect 383 307 385 309
rect 420 308 422 310
rect 430 316 432 318
rect 454 323 456 325
rect 472 323 474 325
rect 495 315 497 317
rect 509 316 511 318
rect 464 307 466 309
rect 483 307 485 309
rect 520 308 522 310
rect 530 316 532 318
rect 554 323 556 325
rect 572 323 574 325
rect 595 315 597 317
rect 609 316 611 318
rect 564 307 566 309
rect 583 307 585 309
rect 620 308 622 310
rect 630 316 632 318
rect 654 323 656 325
rect 672 323 674 325
rect 695 315 697 317
rect 709 316 711 318
rect 664 307 666 309
rect 683 307 685 309
rect 720 308 722 310
rect 730 316 732 318
rect 754 323 756 325
rect 772 323 774 325
rect 795 315 797 317
rect 764 307 766 309
rect 783 307 785 309
rect 21 277 23 279
rect 40 277 42 279
rect 9 269 11 271
rect 32 261 34 263
rect 50 261 52 263
rect 74 268 76 270
rect 84 276 86 278
rect 121 277 123 279
rect 140 277 142 279
rect 95 268 97 270
rect 109 269 111 271
rect 132 261 134 263
rect 150 261 152 263
rect 174 268 176 270
rect 184 276 186 278
rect 221 277 223 279
rect 240 277 242 279
rect 195 268 197 270
rect 209 269 211 271
rect 232 261 234 263
rect 250 261 252 263
rect 274 268 276 270
rect 284 276 286 278
rect 321 277 323 279
rect 340 277 342 279
rect 295 269 297 271
rect 309 269 311 271
rect 332 261 334 263
rect 350 261 352 263
rect 374 268 376 270
rect 384 276 386 278
rect 423 277 425 279
rect 442 277 444 279
rect 395 268 397 270
rect 411 269 413 271
rect 434 261 436 263
rect 452 261 454 263
rect 476 268 478 270
rect 486 276 488 278
rect 523 277 525 279
rect 542 277 544 279
rect 497 269 499 271
rect 511 269 513 271
rect 534 261 536 263
rect 552 261 554 263
rect 576 268 578 270
rect 586 276 588 278
rect 623 277 625 279
rect 642 277 644 279
rect 597 268 599 270
rect 611 269 613 271
rect 634 261 636 263
rect 652 261 654 263
rect 676 268 678 270
rect 686 276 688 278
rect 723 277 725 279
rect 742 277 744 279
rect 697 269 699 271
rect 711 269 713 271
rect 734 261 736 263
rect 752 261 754 263
rect 776 268 778 270
rect 786 276 788 278
rect 797 268 799 270
rect 9 171 11 173
rect 32 179 34 181
rect 21 163 23 165
rect 40 163 42 165
rect 50 179 52 181
rect 74 172 76 174
rect 95 172 97 174
rect 109 171 111 173
rect 84 164 86 166
rect 132 179 134 181
rect 121 163 123 165
rect 140 163 142 165
rect 150 179 152 181
rect 174 172 176 174
rect 195 172 197 174
rect 209 171 211 173
rect 184 164 186 166
rect 232 179 234 181
rect 221 163 223 165
rect 240 163 242 165
rect 250 179 252 181
rect 274 172 276 174
rect 295 172 297 174
rect 309 171 311 173
rect 284 164 286 166
rect 332 179 334 181
rect 321 163 323 165
rect 340 163 342 165
rect 350 179 352 181
rect 374 172 376 174
rect 395 172 397 174
rect 411 171 413 173
rect 384 164 386 166
rect 434 179 436 181
rect 423 163 425 165
rect 442 163 444 165
rect 452 179 454 181
rect 476 172 478 174
rect 497 172 499 174
rect 511 171 513 173
rect 486 164 488 166
rect 534 179 536 181
rect 523 163 525 165
rect 542 163 544 165
rect 552 179 554 181
rect 576 172 578 174
rect 597 172 599 174
rect 611 171 613 173
rect 586 164 588 166
rect 634 179 636 181
rect 623 163 625 165
rect 642 163 644 165
rect 652 179 654 181
rect 676 172 678 174
rect 697 172 699 174
rect 711 171 713 173
rect 686 164 688 166
rect 734 179 736 181
rect 723 163 725 165
rect 742 163 744 165
rect 752 179 754 181
rect 776 172 778 174
rect 797 172 799 174
rect 786 164 788 166
rect 21 133 23 135
rect 40 133 42 135
rect 9 125 11 127
rect 32 117 34 119
rect 50 117 52 119
rect 74 124 76 126
rect 84 132 86 134
rect 121 133 123 135
rect 140 133 142 135
rect 95 124 97 126
rect 109 125 111 127
rect 132 117 134 119
rect 150 117 152 119
rect 174 124 176 126
rect 184 132 186 134
rect 221 133 223 135
rect 240 133 242 135
rect 195 124 197 126
rect 209 125 211 127
rect 232 117 234 119
rect 250 117 252 119
rect 274 124 276 126
rect 284 132 286 134
rect 321 133 323 135
rect 340 133 342 135
rect 295 124 297 126
rect 309 125 311 127
rect 332 117 334 119
rect 350 117 352 119
rect 374 124 376 126
rect 384 132 386 134
rect 423 133 425 135
rect 442 133 444 135
rect 395 124 397 126
rect 411 125 413 127
rect 434 117 436 119
rect 452 117 454 119
rect 476 124 478 126
rect 486 132 488 134
rect 523 133 525 135
rect 542 133 544 135
rect 497 124 499 126
rect 511 125 513 127
rect 534 117 536 119
rect 552 117 554 119
rect 576 124 578 126
rect 586 132 588 134
rect 623 133 625 135
rect 642 133 644 135
rect 597 124 599 126
rect 611 125 613 127
rect 634 117 636 119
rect 652 117 654 119
rect 676 124 678 126
rect 686 132 688 134
rect 723 133 725 135
rect 742 133 744 135
rect 697 124 699 126
rect 711 125 713 127
rect 734 117 736 119
rect 752 117 754 119
rect 776 124 778 126
rect 786 132 788 134
rect 797 124 799 126
rect 9 28 11 30
rect 20 20 22 22
rect 30 28 32 30
rect 54 35 56 37
rect 72 35 74 37
rect 95 27 97 29
rect 64 19 66 21
rect 83 19 85 21
rect 120 20 122 22
rect 130 28 132 30
rect 154 35 156 37
rect 172 35 174 37
rect 195 27 197 29
rect 209 28 211 30
rect 164 19 166 21
rect 183 19 185 21
rect 220 20 222 22
rect 230 28 232 30
rect 254 35 256 37
rect 272 35 274 37
rect 295 27 297 29
rect 309 28 311 30
rect 264 19 266 21
rect 283 19 285 21
rect 320 20 322 22
rect 330 28 332 30
rect 354 35 356 37
rect 372 35 374 37
rect 395 27 397 29
rect 409 28 411 30
rect 364 19 366 21
rect 383 19 385 21
rect 420 20 422 22
rect 430 28 432 30
rect 454 35 456 37
rect 472 35 474 37
rect 495 27 497 29
rect 509 28 511 30
rect 464 19 466 21
rect 483 19 485 21
rect 520 20 522 22
rect 530 28 532 30
rect 554 35 556 37
rect 572 35 574 37
rect 595 27 597 29
rect 609 28 611 30
rect 564 19 566 21
rect 583 19 585 21
rect 620 20 622 22
rect 630 28 632 30
rect 654 35 656 37
rect 672 35 674 37
rect 695 27 697 29
rect 709 28 711 30
rect 664 19 666 21
rect 683 19 685 21
rect 720 20 722 22
rect 730 28 732 30
rect 754 35 756 37
rect 772 35 774 37
rect 795 27 797 29
rect 764 19 766 21
rect 783 19 785 21
<< pdifct1 >>
rect 40 323 42 325
rect 40 316 42 318
rect 40 309 42 311
rect 109 316 111 318
rect 140 323 142 325
rect 140 316 142 318
rect 140 309 142 311
rect 240 323 242 325
rect 240 316 242 318
rect 240 309 242 311
rect 340 316 342 318
rect 340 309 342 311
rect 440 323 442 325
rect 440 316 442 318
rect 440 309 442 311
rect 540 323 542 325
rect 540 316 542 318
rect 540 309 542 311
rect 640 323 642 325
rect 640 316 642 318
rect 640 309 642 311
rect 740 323 742 325
rect 740 316 742 318
rect 740 309 742 311
rect 64 275 66 277
rect 64 268 66 270
rect 64 261 66 263
rect 164 275 166 277
rect 164 268 166 270
rect 164 261 166 263
rect 264 275 266 277
rect 264 268 266 270
rect 264 261 266 263
rect 364 275 366 277
rect 364 268 366 270
rect 364 261 366 263
rect 466 275 468 277
rect 466 268 468 270
rect 466 261 468 263
rect 566 275 568 277
rect 566 268 568 270
rect 566 261 568 263
rect 666 275 668 277
rect 666 268 668 270
rect 666 261 668 263
rect 766 275 768 277
rect 766 268 768 270
rect 766 261 768 263
rect 64 179 66 181
rect 64 172 66 174
rect 64 165 66 167
rect 164 179 166 181
rect 164 172 166 174
rect 164 165 166 167
rect 264 179 266 181
rect 264 172 266 174
rect 264 165 266 167
rect 364 179 366 181
rect 364 172 366 174
rect 364 165 366 167
rect 466 179 468 181
rect 466 172 468 174
rect 466 165 468 167
rect 566 179 568 181
rect 566 172 568 174
rect 566 165 568 167
rect 666 179 668 181
rect 666 172 668 174
rect 666 165 668 167
rect 766 179 768 181
rect 766 172 768 174
rect 766 165 768 167
rect 64 131 66 133
rect 64 124 66 126
rect 64 117 66 119
rect 164 131 166 133
rect 164 124 166 126
rect 164 117 166 119
rect 264 131 266 133
rect 264 124 266 126
rect 264 117 266 119
rect 364 131 366 133
rect 364 124 366 126
rect 364 117 366 119
rect 466 131 468 133
rect 466 124 468 126
rect 466 117 468 119
rect 566 131 568 133
rect 566 124 568 126
rect 566 117 568 119
rect 666 131 668 133
rect 666 124 668 126
rect 666 117 668 119
rect 766 131 768 133
rect 766 124 768 126
rect 766 117 768 119
rect 40 35 42 37
rect 40 28 42 30
rect 40 21 42 23
rect 109 28 111 30
rect 140 35 142 37
rect 140 28 142 30
rect 140 21 142 23
rect 240 35 242 37
rect 240 28 242 30
rect 240 21 242 23
rect 340 35 342 37
rect 340 28 342 30
rect 340 21 342 23
rect 440 35 442 37
rect 440 28 442 30
rect 440 21 442 23
rect 540 35 542 37
rect 540 28 542 30
rect 540 21 542 23
rect 640 35 642 37
rect 640 28 642 30
rect 640 21 642 23
rect 740 35 742 37
rect 740 28 742 30
rect 740 21 742 23
<< alu0 >>
rect 20 349 26 357
rect 61 351 65 357
rect 83 355 84 357
rect 86 355 88 357
rect 83 354 88 355
rect 20 347 22 349
rect 24 347 26 349
rect 20 346 26 347
rect 50 349 57 350
rect 50 347 52 349
rect 54 347 57 349
rect 61 349 62 351
rect 64 349 65 351
rect 61 347 65 349
rect 50 346 57 347
rect 10 344 14 346
rect 10 342 11 344
rect 13 343 14 344
rect 31 344 35 346
rect 13 342 28 343
rect 10 339 28 342
rect 24 334 28 339
rect 24 332 25 334
rect 27 332 28 334
rect 24 327 28 332
rect 20 323 28 327
rect 31 342 32 344
rect 34 342 35 344
rect 20 319 24 323
rect 31 319 35 342
rect 7 318 24 319
rect 7 316 9 318
rect 11 316 24 318
rect 7 315 24 316
rect 28 318 35 319
rect 28 316 30 318
rect 32 316 35 318
rect 28 315 35 316
rect 46 334 50 336
rect 46 332 47 334
rect 49 332 50 334
rect 46 318 50 332
rect 53 325 57 346
rect 69 346 75 348
rect 69 344 72 346
rect 74 344 75 346
rect 69 342 75 344
rect 69 335 73 342
rect 60 334 73 335
rect 60 332 62 334
rect 64 332 73 334
rect 120 349 126 357
rect 161 351 165 357
rect 182 355 184 357
rect 186 355 188 357
rect 182 354 188 355
rect 94 346 99 348
rect 120 347 122 349
rect 124 347 126 349
rect 120 346 126 347
rect 150 349 157 350
rect 150 347 152 349
rect 154 347 157 349
rect 161 349 162 351
rect 164 349 165 351
rect 161 347 165 349
rect 150 346 157 347
rect 94 344 95 346
rect 97 344 99 346
rect 94 342 99 344
rect 60 331 73 332
rect 53 323 54 325
rect 56 323 57 325
rect 53 321 57 323
rect 69 327 73 331
rect 69 325 75 327
rect 69 323 72 325
rect 74 323 75 325
rect 69 321 75 323
rect 95 318 99 342
rect 110 344 114 346
rect 110 342 111 344
rect 113 343 114 344
rect 131 344 135 346
rect 113 342 128 343
rect 110 339 128 342
rect 124 334 128 339
rect 124 332 125 334
rect 127 332 128 334
rect 124 327 128 332
rect 120 323 128 327
rect 131 342 132 344
rect 134 342 135 344
rect 120 319 124 323
rect 131 319 135 342
rect 46 317 99 318
rect 46 315 95 317
rect 97 315 99 317
rect 111 315 124 319
rect 128 318 135 319
rect 128 316 130 318
rect 132 316 135 318
rect 128 315 135 316
rect 46 314 99 315
rect 146 334 150 336
rect 146 332 147 334
rect 149 332 150 334
rect 146 318 150 332
rect 153 325 157 346
rect 169 346 175 348
rect 169 344 172 346
rect 174 344 175 346
rect 169 342 175 344
rect 169 335 173 342
rect 160 334 173 335
rect 160 332 162 334
rect 164 332 173 334
rect 220 349 226 357
rect 261 351 265 357
rect 282 355 284 357
rect 286 355 288 357
rect 282 354 288 355
rect 194 346 199 348
rect 220 347 222 349
rect 224 347 226 349
rect 220 346 226 347
rect 250 349 257 350
rect 250 347 252 349
rect 254 347 257 349
rect 261 349 262 351
rect 264 349 265 351
rect 261 347 265 349
rect 250 346 257 347
rect 194 344 195 346
rect 197 344 199 346
rect 194 342 199 344
rect 160 331 173 332
rect 153 323 154 325
rect 156 323 157 325
rect 153 321 157 323
rect 169 327 173 331
rect 169 325 175 327
rect 169 323 172 325
rect 174 323 175 325
rect 169 321 175 323
rect 195 318 199 342
rect 210 344 214 346
rect 210 342 211 344
rect 213 343 214 344
rect 231 344 235 346
rect 213 342 228 343
rect 210 339 228 342
rect 224 334 228 339
rect 224 332 225 334
rect 227 332 228 334
rect 224 327 228 332
rect 220 323 228 327
rect 231 342 232 344
rect 234 342 235 344
rect 220 319 224 323
rect 231 319 235 342
rect 146 317 199 318
rect 146 315 195 317
rect 197 315 199 317
rect 207 318 224 319
rect 207 316 209 318
rect 211 316 224 318
rect 207 315 224 316
rect 228 318 235 319
rect 228 316 230 318
rect 232 316 235 318
rect 228 315 235 316
rect 146 314 199 315
rect 246 334 250 336
rect 246 332 247 334
rect 249 332 250 334
rect 246 318 250 332
rect 253 325 257 346
rect 269 346 275 348
rect 269 344 272 346
rect 274 344 275 346
rect 269 342 275 344
rect 269 335 273 342
rect 260 334 273 335
rect 260 332 262 334
rect 264 332 273 334
rect 320 349 326 357
rect 361 351 365 357
rect 382 355 384 357
rect 386 355 388 357
rect 382 354 388 355
rect 294 346 299 348
rect 320 347 322 349
rect 324 347 326 349
rect 320 346 326 347
rect 350 349 357 350
rect 350 347 352 349
rect 354 347 357 349
rect 361 349 362 351
rect 364 349 365 351
rect 361 347 365 349
rect 350 346 357 347
rect 294 344 295 346
rect 297 344 299 346
rect 294 342 299 344
rect 260 331 273 332
rect 253 323 254 325
rect 256 323 257 325
rect 253 321 257 323
rect 269 327 273 331
rect 269 325 275 327
rect 269 323 272 325
rect 274 323 275 325
rect 269 321 275 323
rect 295 318 299 342
rect 310 344 314 346
rect 310 342 311 344
rect 313 343 314 344
rect 331 344 335 346
rect 313 342 328 343
rect 310 339 328 342
rect 324 334 328 339
rect 324 332 325 334
rect 327 332 328 334
rect 324 327 328 332
rect 320 323 328 327
rect 331 342 332 344
rect 334 342 335 344
rect 320 319 324 323
rect 331 319 335 342
rect 246 317 299 318
rect 246 315 295 317
rect 297 315 299 317
rect 307 318 324 319
rect 307 316 309 318
rect 311 316 324 318
rect 307 315 324 316
rect 328 318 335 319
rect 328 316 330 318
rect 332 316 335 318
rect 328 315 335 316
rect 246 314 299 315
rect 346 334 350 336
rect 346 332 347 334
rect 349 332 350 334
rect 346 318 350 332
rect 353 325 357 346
rect 369 346 375 348
rect 420 349 426 357
rect 461 351 465 357
rect 482 355 484 357
rect 486 355 488 357
rect 482 354 488 355
rect 369 344 372 346
rect 374 344 375 346
rect 369 342 375 344
rect 369 335 373 342
rect 394 346 399 348
rect 420 347 422 349
rect 424 347 426 349
rect 420 346 426 347
rect 450 349 457 350
rect 450 347 452 349
rect 454 347 457 349
rect 461 349 462 351
rect 464 349 465 351
rect 461 347 465 349
rect 450 346 457 347
rect 394 344 395 346
rect 397 344 399 346
rect 394 342 399 344
rect 360 334 373 335
rect 360 332 362 334
rect 364 332 373 334
rect 360 331 373 332
rect 353 323 354 325
rect 356 323 357 325
rect 353 321 357 323
rect 369 327 373 331
rect 369 325 375 327
rect 369 323 372 325
rect 374 323 375 325
rect 369 321 375 323
rect 395 318 399 342
rect 410 344 414 346
rect 410 342 411 344
rect 413 343 414 344
rect 431 344 435 346
rect 413 342 428 343
rect 410 339 428 342
rect 424 334 428 339
rect 424 332 425 334
rect 427 332 428 334
rect 424 327 428 332
rect 420 323 428 327
rect 431 342 432 344
rect 434 342 435 344
rect 420 319 424 323
rect 431 319 435 342
rect 346 317 399 318
rect 346 315 395 317
rect 397 315 399 317
rect 407 318 424 319
rect 407 316 409 318
rect 411 316 424 318
rect 407 315 424 316
rect 428 318 435 319
rect 428 316 430 318
rect 432 316 435 318
rect 428 315 435 316
rect 346 314 399 315
rect 446 334 450 336
rect 446 332 447 334
rect 449 332 450 334
rect 446 318 450 332
rect 453 325 457 346
rect 469 346 475 348
rect 469 344 472 346
rect 474 344 475 346
rect 469 342 475 344
rect 469 335 473 342
rect 494 346 499 348
rect 494 344 495 346
rect 497 344 499 346
rect 494 342 499 344
rect 460 334 473 335
rect 460 332 462 334
rect 464 332 473 334
rect 460 331 473 332
rect 453 323 454 325
rect 456 323 457 325
rect 453 321 457 323
rect 469 327 473 331
rect 469 325 475 327
rect 469 323 472 325
rect 474 323 475 325
rect 469 321 475 323
rect 495 318 499 342
rect 520 349 526 357
rect 561 351 565 357
rect 582 355 584 357
rect 586 355 588 357
rect 582 354 588 355
rect 520 347 522 349
rect 524 347 526 349
rect 520 346 526 347
rect 550 349 557 350
rect 550 347 552 349
rect 554 347 557 349
rect 561 349 562 351
rect 564 349 565 351
rect 561 347 565 349
rect 550 346 557 347
rect 510 344 514 346
rect 510 342 511 344
rect 513 343 514 344
rect 531 344 535 346
rect 513 342 528 343
rect 510 339 528 342
rect 524 334 528 339
rect 524 332 525 334
rect 527 332 528 334
rect 524 327 528 332
rect 520 323 528 327
rect 531 342 532 344
rect 534 342 535 344
rect 520 319 524 323
rect 531 319 535 342
rect 446 317 499 318
rect 446 315 495 317
rect 497 315 499 317
rect 507 318 524 319
rect 507 316 509 318
rect 511 316 524 318
rect 507 315 524 316
rect 528 318 535 319
rect 528 316 530 318
rect 532 316 535 318
rect 528 315 535 316
rect 446 314 499 315
rect 546 334 550 336
rect 546 332 547 334
rect 549 332 550 334
rect 546 318 550 332
rect 553 325 557 346
rect 569 346 575 348
rect 569 344 572 346
rect 574 344 575 346
rect 569 342 575 344
rect 569 335 573 342
rect 594 346 599 348
rect 594 344 595 346
rect 597 344 599 346
rect 594 342 599 344
rect 560 334 573 335
rect 560 332 562 334
rect 564 332 573 334
rect 560 331 573 332
rect 553 323 554 325
rect 556 323 557 325
rect 553 321 557 323
rect 569 327 573 331
rect 569 325 575 327
rect 569 323 572 325
rect 574 323 575 325
rect 569 321 575 323
rect 595 318 599 342
rect 620 349 626 357
rect 661 351 665 357
rect 682 355 684 357
rect 686 355 688 357
rect 682 354 688 355
rect 620 347 622 349
rect 624 347 626 349
rect 620 346 626 347
rect 650 349 657 350
rect 650 347 652 349
rect 654 347 657 349
rect 661 349 662 351
rect 664 349 665 351
rect 661 347 665 349
rect 650 346 657 347
rect 610 344 614 346
rect 610 342 611 344
rect 613 343 614 344
rect 631 344 635 346
rect 613 342 628 343
rect 610 339 628 342
rect 624 334 628 339
rect 624 332 625 334
rect 627 332 628 334
rect 624 327 628 332
rect 620 323 628 327
rect 631 342 632 344
rect 634 342 635 344
rect 620 319 624 323
rect 631 319 635 342
rect 546 317 599 318
rect 546 315 595 317
rect 597 315 599 317
rect 607 318 624 319
rect 607 316 609 318
rect 611 316 624 318
rect 607 315 624 316
rect 628 318 635 319
rect 628 316 630 318
rect 632 316 635 318
rect 628 315 635 316
rect 546 314 599 315
rect 646 334 650 336
rect 646 332 647 334
rect 649 332 650 334
rect 646 318 650 332
rect 653 325 657 346
rect 669 346 675 348
rect 669 344 672 346
rect 674 344 675 346
rect 669 342 675 344
rect 669 335 673 342
rect 694 346 699 348
rect 694 344 695 346
rect 697 344 699 346
rect 694 342 699 344
rect 660 334 673 335
rect 660 332 662 334
rect 664 332 673 334
rect 660 331 673 332
rect 653 323 654 325
rect 656 323 657 325
rect 653 321 657 323
rect 669 327 673 331
rect 669 325 675 327
rect 669 323 672 325
rect 674 323 675 325
rect 669 321 675 323
rect 695 318 699 342
rect 720 349 726 357
rect 761 351 765 357
rect 782 355 784 357
rect 786 355 788 357
rect 782 354 788 355
rect 720 347 722 349
rect 724 347 726 349
rect 720 346 726 347
rect 750 349 757 350
rect 750 347 752 349
rect 754 347 757 349
rect 761 349 762 351
rect 764 349 765 351
rect 761 347 765 349
rect 750 346 757 347
rect 710 344 714 346
rect 710 342 711 344
rect 713 343 714 344
rect 731 344 735 346
rect 713 342 728 343
rect 710 339 728 342
rect 724 334 728 339
rect 724 332 725 334
rect 727 332 728 334
rect 724 327 728 332
rect 720 323 728 327
rect 731 342 732 344
rect 734 342 735 344
rect 720 319 724 323
rect 731 319 735 342
rect 646 317 699 318
rect 646 315 695 317
rect 697 315 699 317
rect 707 318 724 319
rect 707 316 709 318
rect 711 316 724 318
rect 707 315 724 316
rect 728 318 735 319
rect 728 316 730 318
rect 732 316 735 318
rect 728 315 735 316
rect 646 314 699 315
rect 746 334 750 336
rect 746 332 747 334
rect 749 332 750 334
rect 746 318 750 332
rect 753 325 757 346
rect 769 346 775 348
rect 769 344 772 346
rect 774 344 775 346
rect 769 342 775 344
rect 769 335 773 342
rect 794 346 799 348
rect 794 344 795 346
rect 797 344 799 346
rect 794 342 799 344
rect 760 334 773 335
rect 760 332 762 334
rect 764 332 773 334
rect 760 331 773 332
rect 753 323 754 325
rect 756 323 757 325
rect 753 321 757 323
rect 769 327 773 331
rect 769 325 775 327
rect 769 323 772 325
rect 774 323 775 325
rect 769 321 775 323
rect 795 318 799 342
rect 746 317 799 318
rect 746 315 795 317
rect 797 315 799 317
rect 746 314 799 315
rect 18 310 24 311
rect 18 308 20 310
rect 22 308 24 310
rect 18 301 24 308
rect 118 310 124 311
rect 62 309 68 310
rect 62 307 64 309
rect 66 307 68 309
rect 62 301 68 307
rect 81 309 87 310
rect 81 307 83 309
rect 85 307 87 309
rect 81 301 87 307
rect 118 308 120 310
rect 122 308 124 310
rect 118 301 124 308
rect 218 310 224 311
rect 162 309 168 310
rect 162 307 164 309
rect 166 307 168 309
rect 162 301 168 307
rect 181 309 187 310
rect 181 307 183 309
rect 185 307 187 309
rect 181 301 187 307
rect 218 308 220 310
rect 222 308 224 310
rect 218 301 224 308
rect 318 310 324 311
rect 262 309 268 310
rect 262 307 264 309
rect 266 307 268 309
rect 262 301 268 307
rect 281 309 287 310
rect 281 307 283 309
rect 285 307 287 309
rect 281 301 287 307
rect 318 308 320 310
rect 322 308 324 310
rect 318 301 324 308
rect 418 310 424 311
rect 362 309 368 310
rect 362 307 364 309
rect 366 307 368 309
rect 362 301 368 307
rect 381 309 387 310
rect 381 307 383 309
rect 385 307 387 309
rect 381 301 387 307
rect 418 308 420 310
rect 422 308 424 310
rect 418 301 424 308
rect 518 310 524 311
rect 462 309 468 310
rect 462 307 464 309
rect 466 307 468 309
rect 462 301 468 307
rect 481 309 487 310
rect 481 307 483 309
rect 485 307 487 309
rect 481 301 487 307
rect 518 308 520 310
rect 522 308 524 310
rect 518 301 524 308
rect 618 310 624 311
rect 562 309 568 310
rect 562 307 564 309
rect 566 307 568 309
rect 562 301 568 307
rect 581 309 587 310
rect 581 307 583 309
rect 585 307 587 309
rect 581 301 587 307
rect 618 308 620 310
rect 622 308 624 310
rect 618 301 624 308
rect 718 310 724 311
rect 662 309 668 310
rect 662 307 664 309
rect 666 307 668 309
rect 662 301 668 307
rect 681 309 687 310
rect 681 307 683 309
rect 685 307 687 309
rect 681 301 687 307
rect 718 308 720 310
rect 722 308 724 310
rect 718 301 724 308
rect 762 309 768 310
rect 762 307 764 309
rect 766 307 768 309
rect 762 301 768 307
rect 781 309 787 310
rect 781 307 783 309
rect 785 307 787 309
rect 781 301 787 307
rect 19 279 25 285
rect 19 277 21 279
rect 23 277 25 279
rect 19 276 25 277
rect 38 279 44 285
rect 38 277 40 279
rect 42 277 44 279
rect 38 276 44 277
rect 82 278 88 285
rect 82 276 84 278
rect 86 276 88 278
rect 119 279 125 285
rect 119 277 121 279
rect 123 277 125 279
rect 119 276 125 277
rect 138 279 144 285
rect 138 277 140 279
rect 142 277 144 279
rect 138 276 144 277
rect 82 275 88 276
rect 182 278 188 285
rect 182 276 184 278
rect 186 276 188 278
rect 219 279 225 285
rect 219 277 221 279
rect 223 277 225 279
rect 219 276 225 277
rect 238 279 244 285
rect 238 277 240 279
rect 242 277 244 279
rect 238 276 244 277
rect 182 275 188 276
rect 282 278 288 285
rect 282 276 284 278
rect 286 276 288 278
rect 319 279 325 285
rect 319 277 321 279
rect 323 277 325 279
rect 319 276 325 277
rect 338 279 344 285
rect 338 277 340 279
rect 342 277 344 279
rect 338 276 344 277
rect 282 275 288 276
rect 382 278 388 285
rect 382 276 384 278
rect 386 276 388 278
rect 421 279 427 285
rect 421 277 423 279
rect 425 277 427 279
rect 421 276 427 277
rect 440 279 446 285
rect 440 277 442 279
rect 444 277 446 279
rect 440 276 446 277
rect 382 275 388 276
rect 484 278 490 285
rect 484 276 486 278
rect 488 276 490 278
rect 521 279 527 285
rect 521 277 523 279
rect 525 277 527 279
rect 521 276 527 277
rect 540 279 546 285
rect 540 277 542 279
rect 544 277 546 279
rect 540 276 546 277
rect 484 275 490 276
rect 584 278 590 285
rect 584 276 586 278
rect 588 276 590 278
rect 621 279 627 285
rect 621 277 623 279
rect 625 277 627 279
rect 621 276 627 277
rect 640 279 646 285
rect 640 277 642 279
rect 644 277 646 279
rect 640 276 646 277
rect 584 275 590 276
rect 684 278 690 285
rect 684 276 686 278
rect 688 276 690 278
rect 721 279 727 285
rect 721 277 723 279
rect 725 277 727 279
rect 721 276 727 277
rect 740 279 746 285
rect 740 277 742 279
rect 744 277 746 279
rect 740 276 746 277
rect 684 275 690 276
rect 784 278 790 285
rect 784 276 786 278
rect 788 276 790 278
rect 784 275 790 276
rect 7 271 60 272
rect 7 269 9 271
rect 11 269 60 271
rect 7 268 60 269
rect 7 244 11 268
rect 31 263 37 265
rect 31 261 32 263
rect 34 261 37 263
rect 31 259 37 261
rect 33 255 37 259
rect 49 263 53 265
rect 49 261 50 263
rect 52 261 53 263
rect 33 254 46 255
rect 33 252 42 254
rect 44 252 46 254
rect 33 251 46 252
rect 7 242 12 244
rect 7 240 9 242
rect 11 240 12 242
rect 7 238 12 240
rect 33 244 37 251
rect 31 242 37 244
rect 31 240 32 242
rect 34 240 37 242
rect 31 238 37 240
rect 49 240 53 261
rect 56 254 60 268
rect 56 252 57 254
rect 59 252 60 254
rect 56 250 60 252
rect 107 271 160 272
rect 71 270 78 271
rect 71 268 74 270
rect 76 268 78 270
rect 71 267 78 268
rect 82 270 98 271
rect 82 268 95 270
rect 97 268 98 270
rect 82 267 98 268
rect 107 269 109 271
rect 111 269 160 271
rect 107 268 160 269
rect 71 244 75 267
rect 82 263 86 267
rect 71 242 72 244
rect 74 242 75 244
rect 78 259 86 263
rect 78 254 82 259
rect 78 252 79 254
rect 81 252 82 254
rect 78 247 82 252
rect 78 244 96 247
rect 78 243 93 244
rect 71 240 75 242
rect 92 242 93 243
rect 95 242 96 244
rect 92 240 96 242
rect 49 239 56 240
rect 41 237 45 239
rect 41 235 42 237
rect 44 235 45 237
rect 49 237 52 239
rect 54 237 56 239
rect 49 236 56 237
rect 80 239 86 240
rect 80 237 82 239
rect 84 237 86 239
rect 18 231 24 232
rect 18 229 20 231
rect 22 229 24 231
rect 41 229 45 235
rect 80 229 86 237
rect 107 244 111 268
rect 131 263 137 265
rect 131 261 132 263
rect 134 261 137 263
rect 131 259 137 261
rect 133 255 137 259
rect 149 263 153 265
rect 149 261 150 263
rect 152 261 153 263
rect 133 254 146 255
rect 133 252 142 254
rect 144 252 146 254
rect 133 251 146 252
rect 107 242 112 244
rect 107 240 109 242
rect 111 240 112 242
rect 107 238 112 240
rect 133 244 137 251
rect 131 242 137 244
rect 131 240 132 242
rect 134 240 137 242
rect 131 238 137 240
rect 149 240 153 261
rect 156 254 160 268
rect 156 252 157 254
rect 159 252 160 254
rect 156 250 160 252
rect 207 271 260 272
rect 171 270 178 271
rect 171 268 174 270
rect 176 268 178 270
rect 171 267 178 268
rect 182 270 199 271
rect 182 268 195 270
rect 197 268 199 270
rect 182 267 199 268
rect 207 269 209 271
rect 211 269 260 271
rect 207 268 260 269
rect 171 244 175 267
rect 182 263 186 267
rect 171 242 172 244
rect 174 242 175 244
rect 178 259 186 263
rect 178 254 182 259
rect 178 252 179 254
rect 181 252 182 254
rect 178 247 182 252
rect 178 244 196 247
rect 178 243 193 244
rect 171 240 175 242
rect 192 242 193 243
rect 195 242 196 244
rect 192 240 196 242
rect 207 244 211 268
rect 231 263 237 265
rect 231 261 232 263
rect 234 261 237 263
rect 231 259 237 261
rect 233 255 237 259
rect 249 263 253 265
rect 249 261 250 263
rect 252 261 253 263
rect 233 254 246 255
rect 233 252 242 254
rect 244 252 246 254
rect 233 251 246 252
rect 207 242 212 244
rect 207 240 209 242
rect 211 240 212 242
rect 149 239 156 240
rect 141 237 145 239
rect 141 235 142 237
rect 144 235 145 237
rect 149 237 152 239
rect 154 237 156 239
rect 149 236 156 237
rect 180 239 186 240
rect 180 237 182 239
rect 184 237 186 239
rect 207 238 212 240
rect 233 244 237 251
rect 231 242 237 244
rect 231 240 232 242
rect 234 240 237 242
rect 118 231 124 232
rect 118 229 120 231
rect 122 229 124 231
rect 141 229 145 235
rect 180 229 186 237
rect 231 238 237 240
rect 249 240 253 261
rect 256 254 260 268
rect 256 252 257 254
rect 259 252 260 254
rect 256 250 260 252
rect 282 271 299 272
rect 271 270 278 271
rect 271 268 274 270
rect 276 268 278 270
rect 271 267 278 268
rect 282 269 295 271
rect 297 269 299 271
rect 282 268 299 269
rect 307 271 360 272
rect 307 269 309 271
rect 311 269 360 271
rect 307 268 360 269
rect 271 244 275 267
rect 282 263 286 268
rect 271 242 272 244
rect 274 242 275 244
rect 278 259 286 263
rect 278 254 282 259
rect 278 252 279 254
rect 281 252 282 254
rect 278 247 282 252
rect 278 244 296 247
rect 278 243 293 244
rect 271 240 275 242
rect 292 242 293 243
rect 295 242 296 244
rect 292 240 296 242
rect 307 244 311 268
rect 331 263 337 265
rect 331 261 332 263
rect 334 261 337 263
rect 331 259 337 261
rect 333 255 337 259
rect 349 263 353 265
rect 349 261 350 263
rect 352 261 353 263
rect 333 254 346 255
rect 333 252 342 254
rect 344 252 346 254
rect 333 251 346 252
rect 307 242 312 244
rect 307 240 309 242
rect 311 240 312 242
rect 249 239 256 240
rect 241 237 245 239
rect 241 235 242 237
rect 244 235 245 237
rect 249 237 252 239
rect 254 237 256 239
rect 249 236 256 237
rect 280 239 286 240
rect 280 237 282 239
rect 284 237 286 239
rect 307 238 312 240
rect 333 244 337 251
rect 331 242 337 244
rect 331 240 332 242
rect 334 240 337 242
rect 218 231 224 232
rect 218 229 220 231
rect 222 229 224 231
rect 241 229 245 235
rect 280 229 286 237
rect 331 238 337 240
rect 349 240 353 261
rect 356 254 360 268
rect 356 252 357 254
rect 359 252 360 254
rect 356 250 360 252
rect 409 271 462 272
rect 371 270 378 271
rect 371 268 374 270
rect 376 268 378 270
rect 371 267 378 268
rect 382 270 399 271
rect 382 268 395 270
rect 397 268 399 270
rect 382 267 399 268
rect 409 269 411 271
rect 413 269 462 271
rect 409 268 462 269
rect 371 244 375 267
rect 382 263 386 267
rect 371 242 372 244
rect 374 242 375 244
rect 378 259 386 263
rect 378 254 382 259
rect 378 252 379 254
rect 381 252 382 254
rect 378 247 382 252
rect 378 244 396 247
rect 378 243 393 244
rect 371 240 375 242
rect 392 242 393 243
rect 395 242 396 244
rect 392 240 396 242
rect 349 239 356 240
rect 341 237 345 239
rect 341 235 342 237
rect 344 235 345 237
rect 349 237 352 239
rect 354 237 356 239
rect 349 236 356 237
rect 380 239 386 240
rect 380 237 382 239
rect 384 237 386 239
rect 318 231 324 232
rect 318 229 320 231
rect 322 229 324 231
rect 341 229 345 235
rect 380 229 386 237
rect 409 244 413 268
rect 433 263 439 265
rect 433 261 434 263
rect 436 261 439 263
rect 433 259 439 261
rect 435 255 439 259
rect 451 263 455 265
rect 451 261 452 263
rect 454 261 455 263
rect 435 254 448 255
rect 435 252 444 254
rect 446 252 448 254
rect 435 251 448 252
rect 409 242 414 244
rect 409 240 411 242
rect 413 240 414 242
rect 409 238 414 240
rect 435 244 439 251
rect 433 242 439 244
rect 433 240 434 242
rect 436 240 439 242
rect 433 238 439 240
rect 451 240 455 261
rect 458 254 462 268
rect 458 252 459 254
rect 461 252 462 254
rect 458 250 462 252
rect 484 271 501 272
rect 473 270 480 271
rect 473 268 476 270
rect 478 268 480 270
rect 473 267 480 268
rect 484 269 497 271
rect 499 269 501 271
rect 484 268 501 269
rect 509 271 562 272
rect 509 269 511 271
rect 513 269 562 271
rect 509 268 562 269
rect 473 244 477 267
rect 484 263 488 268
rect 473 242 474 244
rect 476 242 477 244
rect 480 259 488 263
rect 480 254 484 259
rect 480 252 481 254
rect 483 252 484 254
rect 480 247 484 252
rect 480 244 498 247
rect 480 243 495 244
rect 473 240 477 242
rect 494 242 495 243
rect 497 242 498 244
rect 494 240 498 242
rect 509 244 513 268
rect 533 263 539 265
rect 533 261 534 263
rect 536 261 539 263
rect 533 259 539 261
rect 535 255 539 259
rect 551 263 555 265
rect 551 261 552 263
rect 554 261 555 263
rect 535 254 548 255
rect 535 252 544 254
rect 546 252 548 254
rect 535 251 548 252
rect 509 242 514 244
rect 509 240 511 242
rect 513 240 514 242
rect 451 239 458 240
rect 443 237 447 239
rect 443 235 444 237
rect 446 235 447 237
rect 451 237 454 239
rect 456 237 458 239
rect 451 236 458 237
rect 482 239 488 240
rect 482 237 484 239
rect 486 237 488 239
rect 509 238 514 240
rect 535 244 539 251
rect 533 242 539 244
rect 533 240 534 242
rect 536 240 539 242
rect 420 231 426 232
rect 420 229 422 231
rect 424 229 426 231
rect 443 229 447 235
rect 482 229 488 237
rect 533 238 539 240
rect 551 240 555 261
rect 558 254 562 268
rect 558 252 559 254
rect 561 252 562 254
rect 558 250 562 252
rect 609 271 662 272
rect 573 270 580 271
rect 573 268 576 270
rect 578 268 580 270
rect 573 267 580 268
rect 584 270 601 271
rect 584 268 597 270
rect 599 268 601 270
rect 584 267 601 268
rect 609 269 611 271
rect 613 269 662 271
rect 609 268 662 269
rect 573 244 577 267
rect 584 263 588 267
rect 573 242 574 244
rect 576 242 577 244
rect 580 259 588 263
rect 580 254 584 259
rect 580 252 581 254
rect 583 252 584 254
rect 580 247 584 252
rect 580 244 598 247
rect 580 243 595 244
rect 573 240 577 242
rect 594 242 595 243
rect 597 242 598 244
rect 594 240 598 242
rect 609 244 613 268
rect 633 263 639 265
rect 633 261 634 263
rect 636 261 639 263
rect 633 259 639 261
rect 635 255 639 259
rect 651 263 655 265
rect 651 261 652 263
rect 654 261 655 263
rect 635 254 648 255
rect 635 252 644 254
rect 646 252 648 254
rect 635 251 648 252
rect 609 242 614 244
rect 609 240 611 242
rect 613 240 614 242
rect 551 239 558 240
rect 543 237 547 239
rect 543 235 544 237
rect 546 235 547 237
rect 551 237 554 239
rect 556 237 558 239
rect 551 236 558 237
rect 582 239 588 240
rect 582 237 584 239
rect 586 237 588 239
rect 609 238 614 240
rect 635 244 639 251
rect 633 242 639 244
rect 633 240 634 242
rect 636 240 639 242
rect 520 231 526 232
rect 520 229 522 231
rect 524 229 526 231
rect 543 229 547 235
rect 582 229 588 237
rect 633 238 639 240
rect 651 240 655 261
rect 658 254 662 268
rect 658 252 659 254
rect 661 252 662 254
rect 658 250 662 252
rect 684 271 701 272
rect 673 270 680 271
rect 673 268 676 270
rect 678 268 680 270
rect 673 267 680 268
rect 684 269 697 271
rect 699 269 701 271
rect 684 268 701 269
rect 709 271 762 272
rect 709 269 711 271
rect 713 269 762 271
rect 709 268 762 269
rect 673 244 677 267
rect 684 263 688 268
rect 673 242 674 244
rect 676 242 677 244
rect 680 259 688 263
rect 680 254 684 259
rect 680 252 681 254
rect 683 252 684 254
rect 680 247 684 252
rect 680 244 698 247
rect 680 243 695 244
rect 673 240 677 242
rect 694 242 695 243
rect 697 242 698 244
rect 694 240 698 242
rect 709 244 713 268
rect 733 263 739 265
rect 733 261 734 263
rect 736 261 739 263
rect 733 259 739 261
rect 735 255 739 259
rect 751 263 755 265
rect 751 261 752 263
rect 754 261 755 263
rect 735 254 748 255
rect 735 252 744 254
rect 746 252 748 254
rect 735 251 748 252
rect 709 242 714 244
rect 709 240 711 242
rect 713 240 714 242
rect 651 239 658 240
rect 643 237 647 239
rect 643 235 644 237
rect 646 235 647 237
rect 651 237 654 239
rect 656 237 658 239
rect 651 236 658 237
rect 682 239 688 240
rect 682 237 684 239
rect 686 237 688 239
rect 709 238 714 240
rect 735 244 739 251
rect 733 242 739 244
rect 733 240 734 242
rect 736 240 739 242
rect 620 231 626 232
rect 620 229 622 231
rect 624 229 626 231
rect 643 229 647 235
rect 682 229 688 237
rect 733 238 739 240
rect 751 240 755 261
rect 758 254 762 268
rect 758 252 759 254
rect 761 252 762 254
rect 758 250 762 252
rect 773 270 780 271
rect 773 268 776 270
rect 778 268 780 270
rect 773 267 780 268
rect 784 270 801 271
rect 784 268 797 270
rect 799 268 801 270
rect 784 267 801 268
rect 773 244 777 267
rect 784 263 788 267
rect 773 242 774 244
rect 776 242 777 244
rect 780 259 788 263
rect 780 254 784 259
rect 780 252 781 254
rect 783 252 784 254
rect 780 247 784 252
rect 780 244 798 247
rect 780 243 795 244
rect 773 240 777 242
rect 794 242 795 243
rect 797 242 798 244
rect 794 240 798 242
rect 751 239 758 240
rect 743 237 747 239
rect 743 235 744 237
rect 746 235 747 237
rect 751 237 754 239
rect 756 237 758 239
rect 751 236 758 237
rect 782 239 788 240
rect 782 237 784 239
rect 786 237 788 239
rect 720 231 726 232
rect 720 229 722 231
rect 724 229 726 231
rect 743 229 747 235
rect 782 229 788 237
rect 18 211 20 213
rect 22 211 24 213
rect 18 210 24 211
rect 41 207 45 213
rect 7 202 12 204
rect 7 200 9 202
rect 11 200 12 202
rect 7 198 12 200
rect 41 205 42 207
rect 44 205 45 207
rect 7 174 11 198
rect 31 202 37 204
rect 41 203 45 205
rect 49 205 56 206
rect 49 203 52 205
rect 54 203 56 205
rect 31 200 32 202
rect 34 200 37 202
rect 31 198 37 200
rect 33 191 37 198
rect 49 202 56 203
rect 80 205 86 213
rect 118 211 120 213
rect 122 211 124 213
rect 118 210 124 211
rect 141 207 145 213
rect 80 203 82 205
rect 84 203 86 205
rect 80 202 86 203
rect 33 190 46 191
rect 33 188 42 190
rect 44 188 46 190
rect 33 187 46 188
rect 33 183 37 187
rect 31 181 37 183
rect 31 179 32 181
rect 34 179 37 181
rect 31 177 37 179
rect 49 181 53 202
rect 49 179 50 181
rect 52 179 53 181
rect 49 177 53 179
rect 56 190 60 192
rect 56 188 57 190
rect 59 188 60 190
rect 56 174 60 188
rect 7 173 60 174
rect 7 171 9 173
rect 11 171 60 173
rect 7 170 60 171
rect 71 200 75 202
rect 71 198 72 200
rect 74 198 75 200
rect 92 200 96 202
rect 92 199 93 200
rect 71 175 75 198
rect 78 198 93 199
rect 95 198 96 200
rect 78 195 96 198
rect 78 190 82 195
rect 78 188 79 190
rect 81 188 82 190
rect 78 183 82 188
rect 107 202 112 204
rect 107 200 109 202
rect 111 200 112 202
rect 107 198 112 200
rect 141 205 142 207
rect 144 205 145 207
rect 78 179 86 183
rect 82 175 86 179
rect 71 174 78 175
rect 71 172 74 174
rect 76 172 78 174
rect 71 171 78 172
rect 82 174 99 175
rect 82 172 95 174
rect 97 172 99 174
rect 82 171 99 172
rect 107 174 111 198
rect 131 202 137 204
rect 141 203 145 205
rect 149 205 156 206
rect 149 203 152 205
rect 154 203 156 205
rect 131 200 132 202
rect 134 200 137 202
rect 131 198 137 200
rect 133 191 137 198
rect 149 202 156 203
rect 180 205 186 213
rect 218 211 220 213
rect 222 211 224 213
rect 218 210 224 211
rect 241 207 245 213
rect 180 203 182 205
rect 184 203 186 205
rect 180 202 186 203
rect 207 202 212 204
rect 133 190 146 191
rect 133 188 142 190
rect 144 188 146 190
rect 133 187 146 188
rect 133 183 137 187
rect 131 181 137 183
rect 131 179 132 181
rect 134 179 137 181
rect 131 177 137 179
rect 149 181 153 202
rect 149 179 150 181
rect 152 179 153 181
rect 149 177 153 179
rect 156 190 160 192
rect 156 188 157 190
rect 159 188 160 190
rect 156 174 160 188
rect 107 173 160 174
rect 107 171 109 173
rect 111 171 160 173
rect 107 170 160 171
rect 171 200 175 202
rect 171 198 172 200
rect 174 198 175 200
rect 192 200 196 202
rect 192 199 193 200
rect 171 175 175 198
rect 178 198 193 199
rect 195 198 196 200
rect 178 195 196 198
rect 207 200 209 202
rect 211 200 212 202
rect 207 198 212 200
rect 241 205 242 207
rect 244 205 245 207
rect 178 190 182 195
rect 178 188 179 190
rect 181 188 182 190
rect 178 183 182 188
rect 178 179 186 183
rect 182 175 186 179
rect 171 174 178 175
rect 171 172 174 174
rect 176 172 178 174
rect 171 171 178 172
rect 182 174 199 175
rect 182 172 195 174
rect 197 172 199 174
rect 182 171 199 172
rect 207 174 211 198
rect 231 202 237 204
rect 241 203 245 205
rect 249 205 256 206
rect 249 203 252 205
rect 254 203 256 205
rect 231 200 232 202
rect 234 200 237 202
rect 231 198 237 200
rect 233 191 237 198
rect 249 202 256 203
rect 280 205 286 213
rect 318 211 320 213
rect 322 211 324 213
rect 318 210 324 211
rect 341 207 345 213
rect 280 203 282 205
rect 284 203 286 205
rect 280 202 286 203
rect 233 190 246 191
rect 233 188 242 190
rect 244 188 246 190
rect 233 187 246 188
rect 233 183 237 187
rect 231 181 237 183
rect 231 179 232 181
rect 234 179 237 181
rect 231 177 237 179
rect 249 181 253 202
rect 249 179 250 181
rect 252 179 253 181
rect 249 177 253 179
rect 256 190 260 192
rect 256 188 257 190
rect 259 188 260 190
rect 256 174 260 188
rect 207 173 260 174
rect 207 171 209 173
rect 211 171 260 173
rect 207 170 260 171
rect 271 200 275 202
rect 271 198 272 200
rect 274 198 275 200
rect 292 200 296 202
rect 292 199 293 200
rect 271 175 275 198
rect 278 198 293 199
rect 295 198 296 200
rect 278 195 296 198
rect 278 190 282 195
rect 278 188 279 190
rect 281 188 282 190
rect 278 183 282 188
rect 307 202 312 204
rect 307 200 309 202
rect 311 200 312 202
rect 307 198 312 200
rect 341 205 342 207
rect 344 205 345 207
rect 278 179 286 183
rect 282 175 286 179
rect 271 174 278 175
rect 271 172 274 174
rect 276 172 278 174
rect 271 171 278 172
rect 282 174 299 175
rect 282 172 295 174
rect 297 172 299 174
rect 282 171 299 172
rect 307 174 311 198
rect 331 202 337 204
rect 341 203 345 205
rect 349 205 356 206
rect 349 203 352 205
rect 354 203 356 205
rect 331 200 332 202
rect 334 200 337 202
rect 331 198 337 200
rect 333 191 337 198
rect 349 202 356 203
rect 380 205 386 213
rect 420 211 422 213
rect 424 211 426 213
rect 420 210 426 211
rect 443 207 447 213
rect 380 203 382 205
rect 384 203 386 205
rect 380 202 386 203
rect 333 190 346 191
rect 333 188 342 190
rect 344 188 346 190
rect 333 187 346 188
rect 333 183 337 187
rect 331 181 337 183
rect 331 179 332 181
rect 334 179 337 181
rect 331 177 337 179
rect 349 181 353 202
rect 349 179 350 181
rect 352 179 353 181
rect 349 177 353 179
rect 356 190 360 192
rect 356 188 357 190
rect 359 188 360 190
rect 356 174 360 188
rect 307 173 360 174
rect 307 171 309 173
rect 311 171 360 173
rect 307 170 360 171
rect 371 200 375 202
rect 371 198 372 200
rect 374 198 375 200
rect 392 200 396 202
rect 392 199 393 200
rect 371 175 375 198
rect 378 198 393 199
rect 395 198 396 200
rect 378 195 396 198
rect 378 190 382 195
rect 378 188 379 190
rect 381 188 382 190
rect 378 183 382 188
rect 409 202 414 204
rect 409 200 411 202
rect 413 200 414 202
rect 409 198 414 200
rect 443 205 444 207
rect 446 205 447 207
rect 378 179 386 183
rect 382 175 386 179
rect 371 174 378 175
rect 371 172 374 174
rect 376 172 378 174
rect 371 171 378 172
rect 382 174 399 175
rect 382 172 395 174
rect 397 172 399 174
rect 382 171 399 172
rect 409 174 413 198
rect 433 202 439 204
rect 443 203 447 205
rect 451 205 458 206
rect 451 203 454 205
rect 456 203 458 205
rect 433 200 434 202
rect 436 200 439 202
rect 433 198 439 200
rect 435 191 439 198
rect 451 202 458 203
rect 482 205 488 213
rect 520 211 522 213
rect 524 211 526 213
rect 520 210 526 211
rect 543 207 547 213
rect 482 203 484 205
rect 486 203 488 205
rect 482 202 488 203
rect 509 202 514 204
rect 435 190 448 191
rect 435 188 444 190
rect 446 188 448 190
rect 435 187 448 188
rect 435 183 439 187
rect 433 181 439 183
rect 433 179 434 181
rect 436 179 439 181
rect 433 177 439 179
rect 451 181 455 202
rect 451 179 452 181
rect 454 179 455 181
rect 451 177 455 179
rect 458 190 462 192
rect 458 188 459 190
rect 461 188 462 190
rect 458 174 462 188
rect 409 173 462 174
rect 409 171 411 173
rect 413 171 462 173
rect 409 170 462 171
rect 473 200 477 202
rect 473 198 474 200
rect 476 198 477 200
rect 494 200 498 202
rect 494 199 495 200
rect 473 175 477 198
rect 480 198 495 199
rect 497 198 498 200
rect 480 195 498 198
rect 509 200 511 202
rect 513 200 514 202
rect 509 198 514 200
rect 543 205 544 207
rect 546 205 547 207
rect 480 190 484 195
rect 480 188 481 190
rect 483 188 484 190
rect 480 183 484 188
rect 480 179 488 183
rect 484 175 488 179
rect 473 174 480 175
rect 473 172 476 174
rect 478 172 480 174
rect 473 171 480 172
rect 484 174 501 175
rect 484 172 497 174
rect 499 172 501 174
rect 484 171 501 172
rect 509 174 513 198
rect 533 202 539 204
rect 543 203 547 205
rect 551 205 558 206
rect 551 203 554 205
rect 556 203 558 205
rect 533 200 534 202
rect 536 200 539 202
rect 533 198 539 200
rect 535 191 539 198
rect 551 202 558 203
rect 582 205 588 213
rect 620 211 622 213
rect 624 211 626 213
rect 620 210 626 211
rect 643 207 647 213
rect 582 203 584 205
rect 586 203 588 205
rect 582 202 588 203
rect 609 202 614 204
rect 535 190 548 191
rect 535 188 544 190
rect 546 188 548 190
rect 535 187 548 188
rect 535 183 539 187
rect 533 181 539 183
rect 533 179 534 181
rect 536 179 539 181
rect 533 177 539 179
rect 551 181 555 202
rect 551 179 552 181
rect 554 179 555 181
rect 551 177 555 179
rect 558 190 562 192
rect 558 188 559 190
rect 561 188 562 190
rect 558 174 562 188
rect 509 173 562 174
rect 509 171 511 173
rect 513 171 562 173
rect 509 170 562 171
rect 573 200 577 202
rect 573 198 574 200
rect 576 198 577 200
rect 594 200 598 202
rect 594 199 595 200
rect 573 175 577 198
rect 580 198 595 199
rect 597 198 598 200
rect 580 195 598 198
rect 609 200 611 202
rect 613 200 614 202
rect 609 198 614 200
rect 643 205 644 207
rect 646 205 647 207
rect 580 190 584 195
rect 580 188 581 190
rect 583 188 584 190
rect 580 183 584 188
rect 580 179 588 183
rect 584 175 588 179
rect 573 174 580 175
rect 573 172 576 174
rect 578 172 580 174
rect 573 171 580 172
rect 584 174 601 175
rect 584 172 597 174
rect 599 172 601 174
rect 584 171 601 172
rect 609 174 613 198
rect 633 202 639 204
rect 643 203 647 205
rect 651 205 658 206
rect 651 203 654 205
rect 656 203 658 205
rect 633 200 634 202
rect 636 200 639 202
rect 633 198 639 200
rect 635 191 639 198
rect 651 202 658 203
rect 682 205 688 213
rect 720 211 722 213
rect 724 211 726 213
rect 720 210 726 211
rect 743 207 747 213
rect 682 203 684 205
rect 686 203 688 205
rect 682 202 688 203
rect 709 202 714 204
rect 635 190 648 191
rect 635 188 644 190
rect 646 188 648 190
rect 635 187 648 188
rect 635 183 639 187
rect 633 181 639 183
rect 633 179 634 181
rect 636 179 639 181
rect 633 177 639 179
rect 651 181 655 202
rect 651 179 652 181
rect 654 179 655 181
rect 651 177 655 179
rect 658 190 662 192
rect 658 188 659 190
rect 661 188 662 190
rect 658 174 662 188
rect 609 173 662 174
rect 609 171 611 173
rect 613 171 662 173
rect 609 170 662 171
rect 673 200 677 202
rect 673 198 674 200
rect 676 198 677 200
rect 694 200 698 202
rect 694 199 695 200
rect 673 175 677 198
rect 680 198 695 199
rect 697 198 698 200
rect 680 195 698 198
rect 709 200 711 202
rect 713 200 714 202
rect 709 198 714 200
rect 743 205 744 207
rect 746 205 747 207
rect 680 190 684 195
rect 680 188 681 190
rect 683 188 684 190
rect 680 183 684 188
rect 680 179 688 183
rect 684 175 688 179
rect 673 174 680 175
rect 673 172 676 174
rect 678 172 680 174
rect 673 171 680 172
rect 684 174 701 175
rect 684 172 697 174
rect 699 172 701 174
rect 684 171 701 172
rect 709 174 713 198
rect 733 202 739 204
rect 743 203 747 205
rect 751 205 758 206
rect 751 203 754 205
rect 756 203 758 205
rect 733 200 734 202
rect 736 200 739 202
rect 733 198 739 200
rect 735 191 739 198
rect 751 202 758 203
rect 782 205 788 213
rect 782 203 784 205
rect 786 203 788 205
rect 782 202 788 203
rect 735 190 748 191
rect 735 188 744 190
rect 746 188 748 190
rect 735 187 748 188
rect 735 183 739 187
rect 733 181 739 183
rect 733 179 734 181
rect 736 179 739 181
rect 733 177 739 179
rect 751 181 755 202
rect 751 179 752 181
rect 754 179 755 181
rect 751 177 755 179
rect 758 190 762 192
rect 758 188 759 190
rect 761 188 762 190
rect 758 174 762 188
rect 709 173 762 174
rect 709 171 711 173
rect 713 171 762 173
rect 709 170 762 171
rect 773 200 777 202
rect 773 198 774 200
rect 776 198 777 200
rect 794 200 798 202
rect 794 199 795 200
rect 773 175 777 198
rect 780 198 795 199
rect 797 198 798 200
rect 780 195 798 198
rect 780 190 784 195
rect 780 188 781 190
rect 783 188 784 190
rect 780 183 784 188
rect 780 179 788 183
rect 784 175 788 179
rect 773 174 780 175
rect 773 172 776 174
rect 778 172 780 174
rect 773 171 780 172
rect 784 174 801 175
rect 784 172 797 174
rect 799 172 801 174
rect 784 171 801 172
rect 19 165 25 166
rect 19 163 21 165
rect 23 163 25 165
rect 19 157 25 163
rect 38 165 44 166
rect 38 163 40 165
rect 42 163 44 165
rect 82 166 88 167
rect 82 164 84 166
rect 86 164 88 166
rect 38 157 44 163
rect 82 157 88 164
rect 119 165 125 166
rect 119 163 121 165
rect 123 163 125 165
rect 119 157 125 163
rect 138 165 144 166
rect 138 163 140 165
rect 142 163 144 165
rect 182 166 188 167
rect 182 164 184 166
rect 186 164 188 166
rect 138 157 144 163
rect 182 157 188 164
rect 219 165 225 166
rect 219 163 221 165
rect 223 163 225 165
rect 219 157 225 163
rect 238 165 244 166
rect 238 163 240 165
rect 242 163 244 165
rect 282 166 288 167
rect 282 164 284 166
rect 286 164 288 166
rect 238 157 244 163
rect 282 157 288 164
rect 319 165 325 166
rect 319 163 321 165
rect 323 163 325 165
rect 319 157 325 163
rect 338 165 344 166
rect 338 163 340 165
rect 342 163 344 165
rect 382 166 388 167
rect 382 164 384 166
rect 386 164 388 166
rect 338 157 344 163
rect 382 157 388 164
rect 421 165 427 166
rect 421 163 423 165
rect 425 163 427 165
rect 421 157 427 163
rect 440 165 446 166
rect 440 163 442 165
rect 444 163 446 165
rect 484 166 490 167
rect 484 164 486 166
rect 488 164 490 166
rect 440 157 446 163
rect 484 157 490 164
rect 521 165 527 166
rect 521 163 523 165
rect 525 163 527 165
rect 521 157 527 163
rect 540 165 546 166
rect 540 163 542 165
rect 544 163 546 165
rect 584 166 590 167
rect 584 164 586 166
rect 588 164 590 166
rect 540 157 546 163
rect 584 157 590 164
rect 621 165 627 166
rect 621 163 623 165
rect 625 163 627 165
rect 621 157 627 163
rect 640 165 646 166
rect 640 163 642 165
rect 644 163 646 165
rect 684 166 690 167
rect 684 164 686 166
rect 688 164 690 166
rect 640 157 646 163
rect 684 157 690 164
rect 721 165 727 166
rect 721 163 723 165
rect 725 163 727 165
rect 721 157 727 163
rect 740 165 746 166
rect 740 163 742 165
rect 744 163 746 165
rect 784 166 790 167
rect 784 164 786 166
rect 788 164 790 166
rect 740 157 746 163
rect 784 157 790 164
rect 19 135 25 141
rect 19 133 21 135
rect 23 133 25 135
rect 19 132 25 133
rect 38 135 44 141
rect 38 133 40 135
rect 42 133 44 135
rect 38 132 44 133
rect 82 134 88 141
rect 82 132 84 134
rect 86 132 88 134
rect 119 135 125 141
rect 119 133 121 135
rect 123 133 125 135
rect 119 132 125 133
rect 138 135 144 141
rect 138 133 140 135
rect 142 133 144 135
rect 138 132 144 133
rect 82 131 88 132
rect 182 134 188 141
rect 182 132 184 134
rect 186 132 188 134
rect 219 135 225 141
rect 219 133 221 135
rect 223 133 225 135
rect 219 132 225 133
rect 238 135 244 141
rect 238 133 240 135
rect 242 133 244 135
rect 238 132 244 133
rect 182 131 188 132
rect 282 134 288 141
rect 282 132 284 134
rect 286 132 288 134
rect 319 135 325 141
rect 319 133 321 135
rect 323 133 325 135
rect 319 132 325 133
rect 338 135 344 141
rect 338 133 340 135
rect 342 133 344 135
rect 338 132 344 133
rect 282 131 288 132
rect 382 134 388 141
rect 382 132 384 134
rect 386 132 388 134
rect 421 135 427 141
rect 421 133 423 135
rect 425 133 427 135
rect 421 132 427 133
rect 440 135 446 141
rect 440 133 442 135
rect 444 133 446 135
rect 440 132 446 133
rect 382 131 388 132
rect 484 134 490 141
rect 484 132 486 134
rect 488 132 490 134
rect 521 135 527 141
rect 521 133 523 135
rect 525 133 527 135
rect 521 132 527 133
rect 540 135 546 141
rect 540 133 542 135
rect 544 133 546 135
rect 540 132 546 133
rect 484 131 490 132
rect 584 134 590 141
rect 584 132 586 134
rect 588 132 590 134
rect 621 135 627 141
rect 621 133 623 135
rect 625 133 627 135
rect 621 132 627 133
rect 640 135 646 141
rect 640 133 642 135
rect 644 133 646 135
rect 640 132 646 133
rect 584 131 590 132
rect 684 134 690 141
rect 684 132 686 134
rect 688 132 690 134
rect 721 135 727 141
rect 721 133 723 135
rect 725 133 727 135
rect 721 132 727 133
rect 740 135 746 141
rect 740 133 742 135
rect 744 133 746 135
rect 740 132 746 133
rect 684 131 690 132
rect 784 134 790 141
rect 784 132 786 134
rect 788 132 790 134
rect 784 131 790 132
rect 7 127 60 128
rect 7 125 9 127
rect 11 125 60 127
rect 7 124 60 125
rect 7 100 11 124
rect 31 119 37 121
rect 31 117 32 119
rect 34 117 37 119
rect 31 115 37 117
rect 33 111 37 115
rect 49 119 53 121
rect 49 117 50 119
rect 52 117 53 119
rect 33 110 46 111
rect 33 108 42 110
rect 44 108 46 110
rect 33 107 46 108
rect 7 98 12 100
rect 7 96 9 98
rect 11 96 12 98
rect 7 94 12 96
rect 33 100 37 107
rect 31 98 37 100
rect 31 96 32 98
rect 34 96 37 98
rect 31 94 37 96
rect 49 96 53 117
rect 56 110 60 124
rect 56 108 57 110
rect 59 108 60 110
rect 56 106 60 108
rect 107 127 160 128
rect 71 126 78 127
rect 71 124 74 126
rect 76 124 78 126
rect 71 123 78 124
rect 82 126 99 127
rect 82 124 95 126
rect 97 124 99 126
rect 82 123 99 124
rect 107 125 109 127
rect 111 125 160 127
rect 107 124 160 125
rect 71 100 75 123
rect 82 119 86 123
rect 71 98 72 100
rect 74 98 75 100
rect 78 115 86 119
rect 78 110 82 115
rect 78 108 79 110
rect 81 108 82 110
rect 78 103 82 108
rect 78 100 96 103
rect 78 99 93 100
rect 71 96 75 98
rect 92 98 93 99
rect 95 98 96 100
rect 92 96 96 98
rect 107 100 111 124
rect 131 119 137 121
rect 131 117 132 119
rect 134 117 137 119
rect 131 115 137 117
rect 133 111 137 115
rect 149 119 153 121
rect 149 117 150 119
rect 152 117 153 119
rect 133 110 146 111
rect 133 108 142 110
rect 144 108 146 110
rect 133 107 146 108
rect 107 98 112 100
rect 107 96 109 98
rect 111 96 112 98
rect 49 95 56 96
rect 41 93 45 95
rect 41 91 42 93
rect 44 91 45 93
rect 49 93 52 95
rect 54 93 56 95
rect 49 92 56 93
rect 80 95 86 96
rect 80 93 82 95
rect 84 93 86 95
rect 107 94 112 96
rect 133 100 137 107
rect 131 98 137 100
rect 131 96 132 98
rect 134 96 137 98
rect 131 94 137 96
rect 149 96 153 117
rect 156 110 160 124
rect 156 108 157 110
rect 159 108 160 110
rect 156 106 160 108
rect 207 127 260 128
rect 171 126 178 127
rect 171 124 174 126
rect 176 124 178 126
rect 171 123 178 124
rect 182 126 199 127
rect 182 124 195 126
rect 197 124 199 126
rect 182 123 199 124
rect 207 125 209 127
rect 211 125 260 127
rect 207 124 260 125
rect 171 100 175 123
rect 182 119 186 123
rect 171 98 172 100
rect 174 98 175 100
rect 178 115 186 119
rect 178 110 182 115
rect 178 108 179 110
rect 181 108 182 110
rect 178 103 182 108
rect 178 100 196 103
rect 178 99 193 100
rect 171 96 175 98
rect 192 98 193 99
rect 195 98 196 100
rect 192 96 196 98
rect 207 100 211 124
rect 231 119 237 121
rect 231 117 232 119
rect 234 117 237 119
rect 231 115 237 117
rect 233 111 237 115
rect 249 119 253 121
rect 249 117 250 119
rect 252 117 253 119
rect 233 110 246 111
rect 207 98 212 100
rect 207 96 209 98
rect 211 96 212 98
rect 149 95 156 96
rect 18 87 24 88
rect 18 85 20 87
rect 22 85 24 87
rect 41 85 45 91
rect 80 85 86 93
rect 141 93 145 95
rect 141 91 142 93
rect 144 91 145 93
rect 149 93 152 95
rect 154 93 156 95
rect 149 92 156 93
rect 180 95 186 96
rect 180 93 182 95
rect 184 93 186 95
rect 207 94 212 96
rect 233 108 242 110
rect 244 108 246 110
rect 233 107 246 108
rect 233 100 237 107
rect 231 98 237 100
rect 231 96 232 98
rect 234 96 237 98
rect 231 94 237 96
rect 249 96 253 117
rect 256 110 260 124
rect 256 108 257 110
rect 259 108 260 110
rect 256 106 260 108
rect 307 127 360 128
rect 271 126 278 127
rect 271 124 274 126
rect 276 124 278 126
rect 271 123 278 124
rect 282 126 299 127
rect 282 124 295 126
rect 297 124 299 126
rect 282 123 299 124
rect 307 125 309 127
rect 311 125 360 127
rect 307 124 360 125
rect 271 100 275 123
rect 282 119 286 123
rect 271 98 272 100
rect 274 98 275 100
rect 278 115 286 119
rect 278 110 282 115
rect 278 108 279 110
rect 281 108 282 110
rect 278 103 282 108
rect 278 100 296 103
rect 278 99 293 100
rect 271 96 275 98
rect 292 98 293 99
rect 295 98 296 100
rect 292 96 296 98
rect 307 100 311 124
rect 331 119 337 121
rect 331 117 332 119
rect 334 117 337 119
rect 331 115 337 117
rect 333 111 337 115
rect 349 119 353 121
rect 349 117 350 119
rect 352 117 353 119
rect 333 110 346 111
rect 333 108 342 110
rect 344 108 346 110
rect 333 107 346 108
rect 307 98 312 100
rect 307 96 309 98
rect 311 96 312 98
rect 249 95 256 96
rect 118 87 124 88
rect 118 85 120 87
rect 122 85 124 87
rect 141 85 145 91
rect 180 85 186 93
rect 241 93 245 95
rect 241 91 242 93
rect 244 91 245 93
rect 249 93 252 95
rect 254 93 256 95
rect 249 92 256 93
rect 280 95 286 96
rect 280 93 282 95
rect 284 93 286 95
rect 307 94 312 96
rect 333 100 337 107
rect 331 98 337 100
rect 331 96 332 98
rect 334 96 337 98
rect 331 94 337 96
rect 349 96 353 117
rect 356 110 360 124
rect 356 108 357 110
rect 359 108 360 110
rect 356 106 360 108
rect 409 127 462 128
rect 371 126 378 127
rect 371 124 374 126
rect 376 124 378 126
rect 371 123 378 124
rect 382 126 399 127
rect 382 124 395 126
rect 397 124 399 126
rect 382 123 399 124
rect 409 125 411 127
rect 413 125 462 127
rect 409 124 462 125
rect 371 100 375 123
rect 382 119 386 123
rect 371 98 372 100
rect 374 98 375 100
rect 378 115 386 119
rect 378 110 382 115
rect 378 108 379 110
rect 381 108 382 110
rect 378 103 382 108
rect 378 100 396 103
rect 378 99 393 100
rect 371 96 375 98
rect 392 98 393 99
rect 395 98 396 100
rect 392 96 396 98
rect 409 100 413 124
rect 433 119 439 121
rect 433 117 434 119
rect 436 117 439 119
rect 433 115 439 117
rect 435 111 439 115
rect 451 119 455 121
rect 451 117 452 119
rect 454 117 455 119
rect 435 110 448 111
rect 435 108 444 110
rect 446 108 448 110
rect 435 107 448 108
rect 409 98 414 100
rect 409 96 411 98
rect 413 96 414 98
rect 349 95 356 96
rect 218 87 224 88
rect 218 85 220 87
rect 222 85 224 87
rect 241 85 245 91
rect 280 85 286 93
rect 341 93 345 95
rect 341 91 342 93
rect 344 91 345 93
rect 349 93 352 95
rect 354 93 356 95
rect 349 92 356 93
rect 380 95 386 96
rect 380 93 382 95
rect 384 93 386 95
rect 409 94 414 96
rect 435 100 439 107
rect 433 98 439 100
rect 433 96 434 98
rect 436 96 439 98
rect 433 94 439 96
rect 451 96 455 117
rect 458 110 462 124
rect 458 108 459 110
rect 461 108 462 110
rect 458 106 462 108
rect 509 127 562 128
rect 473 126 480 127
rect 473 124 476 126
rect 478 124 480 126
rect 473 123 480 124
rect 484 126 501 127
rect 484 124 497 126
rect 499 124 501 126
rect 484 123 501 124
rect 509 125 511 127
rect 513 125 562 127
rect 509 124 562 125
rect 473 100 477 123
rect 484 119 488 123
rect 473 98 474 100
rect 476 98 477 100
rect 480 115 488 119
rect 480 110 484 115
rect 480 108 481 110
rect 483 108 484 110
rect 480 103 484 108
rect 480 100 498 103
rect 480 99 495 100
rect 473 96 477 98
rect 494 98 495 99
rect 497 98 498 100
rect 494 96 498 98
rect 509 100 513 124
rect 533 119 539 121
rect 533 117 534 119
rect 536 117 539 119
rect 533 115 539 117
rect 535 111 539 115
rect 551 119 555 121
rect 551 117 552 119
rect 554 117 555 119
rect 535 110 548 111
rect 535 108 544 110
rect 546 108 548 110
rect 535 107 548 108
rect 509 98 514 100
rect 509 96 511 98
rect 513 96 514 98
rect 451 95 458 96
rect 318 87 324 88
rect 318 85 320 87
rect 322 85 324 87
rect 341 85 345 91
rect 380 85 386 93
rect 443 93 447 95
rect 443 91 444 93
rect 446 91 447 93
rect 451 93 454 95
rect 456 93 458 95
rect 451 92 458 93
rect 482 95 488 96
rect 482 93 484 95
rect 486 93 488 95
rect 509 94 514 96
rect 535 100 539 107
rect 533 98 539 100
rect 533 96 534 98
rect 536 96 539 98
rect 533 94 539 96
rect 551 96 555 117
rect 558 110 562 124
rect 558 108 559 110
rect 561 108 562 110
rect 558 106 562 108
rect 609 127 662 128
rect 573 126 580 127
rect 573 124 576 126
rect 578 124 580 126
rect 573 123 580 124
rect 584 126 601 127
rect 584 124 597 126
rect 599 124 601 126
rect 584 123 601 124
rect 609 125 611 127
rect 613 125 662 127
rect 609 124 662 125
rect 573 100 577 123
rect 584 119 588 123
rect 573 98 574 100
rect 576 98 577 100
rect 580 115 588 119
rect 580 110 584 115
rect 580 108 581 110
rect 583 108 584 110
rect 580 103 584 108
rect 580 100 598 103
rect 609 100 613 124
rect 633 119 639 121
rect 633 117 634 119
rect 636 117 639 119
rect 633 115 639 117
rect 635 111 639 115
rect 651 119 655 121
rect 651 117 652 119
rect 654 117 655 119
rect 635 110 648 111
rect 635 108 644 110
rect 646 108 648 110
rect 635 107 648 108
rect 580 99 595 100
rect 573 96 577 98
rect 594 98 595 99
rect 597 98 598 100
rect 594 96 598 98
rect 609 98 614 100
rect 609 96 611 98
rect 613 96 614 98
rect 551 95 558 96
rect 420 87 426 88
rect 420 85 422 87
rect 424 85 426 87
rect 443 85 447 91
rect 482 85 488 93
rect 543 93 547 95
rect 543 91 544 93
rect 546 91 547 93
rect 551 93 554 95
rect 556 93 558 95
rect 551 92 558 93
rect 582 95 588 96
rect 582 93 584 95
rect 586 93 588 95
rect 609 94 614 96
rect 635 100 639 107
rect 633 98 639 100
rect 633 96 634 98
rect 636 96 639 98
rect 633 94 639 96
rect 651 96 655 117
rect 658 110 662 124
rect 658 108 659 110
rect 661 108 662 110
rect 658 106 662 108
rect 709 127 762 128
rect 673 126 680 127
rect 673 124 676 126
rect 678 124 680 126
rect 673 123 680 124
rect 684 126 701 127
rect 684 124 697 126
rect 699 124 701 126
rect 684 123 701 124
rect 709 125 711 127
rect 713 125 762 127
rect 709 124 762 125
rect 673 100 677 123
rect 684 119 688 123
rect 673 98 674 100
rect 676 98 677 100
rect 680 115 688 119
rect 680 110 684 115
rect 680 108 681 110
rect 683 108 684 110
rect 680 103 684 108
rect 680 100 698 103
rect 680 99 695 100
rect 673 96 677 98
rect 694 98 695 99
rect 697 98 698 100
rect 694 96 698 98
rect 709 100 713 124
rect 733 119 739 121
rect 733 117 734 119
rect 736 117 739 119
rect 733 115 739 117
rect 735 111 739 115
rect 751 119 755 121
rect 751 117 752 119
rect 754 117 755 119
rect 735 110 748 111
rect 709 98 714 100
rect 709 96 711 98
rect 713 96 714 98
rect 651 95 658 96
rect 520 87 526 88
rect 520 85 522 87
rect 524 85 526 87
rect 543 85 547 91
rect 582 85 588 93
rect 643 93 647 95
rect 643 91 644 93
rect 646 91 647 93
rect 651 93 654 95
rect 656 93 658 95
rect 651 92 658 93
rect 682 95 688 96
rect 682 93 684 95
rect 686 93 688 95
rect 709 94 714 96
rect 735 108 744 110
rect 746 108 748 110
rect 735 107 748 108
rect 735 100 739 107
rect 733 98 739 100
rect 733 96 734 98
rect 736 96 739 98
rect 733 94 739 96
rect 751 96 755 117
rect 758 110 762 124
rect 758 108 759 110
rect 761 108 762 110
rect 758 106 762 108
rect 773 126 780 127
rect 773 124 776 126
rect 778 124 780 126
rect 773 123 780 124
rect 784 126 801 127
rect 784 124 797 126
rect 799 124 801 126
rect 784 123 801 124
rect 773 100 777 123
rect 784 119 788 123
rect 773 98 774 100
rect 776 98 777 100
rect 780 115 788 119
rect 780 110 784 115
rect 780 108 781 110
rect 783 108 784 110
rect 780 103 784 108
rect 780 100 798 103
rect 780 99 795 100
rect 773 96 777 98
rect 794 98 795 99
rect 797 98 798 100
rect 794 96 798 98
rect 751 95 758 96
rect 620 87 626 88
rect 620 85 622 87
rect 624 85 626 87
rect 643 85 647 91
rect 682 85 688 93
rect 743 93 747 95
rect 743 91 744 93
rect 746 91 747 93
rect 751 93 754 95
rect 756 93 758 95
rect 751 92 758 93
rect 782 95 788 96
rect 782 93 784 95
rect 786 93 788 95
rect 720 87 726 88
rect 720 85 722 87
rect 724 85 726 87
rect 743 85 747 91
rect 782 85 788 93
rect 20 61 26 69
rect 61 63 65 69
rect 83 67 84 69
rect 86 67 88 69
rect 83 66 88 67
rect 20 59 22 61
rect 24 59 26 61
rect 20 58 26 59
rect 50 61 57 62
rect 50 59 52 61
rect 54 59 57 61
rect 61 61 62 63
rect 64 61 65 63
rect 61 59 65 61
rect 50 58 57 59
rect 10 56 14 58
rect 10 54 11 56
rect 13 55 14 56
rect 31 56 35 58
rect 13 54 28 55
rect 10 51 28 54
rect 24 46 28 51
rect 24 44 25 46
rect 27 44 28 46
rect 24 39 28 44
rect 20 35 28 39
rect 31 54 32 56
rect 34 54 35 56
rect 20 31 24 35
rect 31 31 35 54
rect 7 30 24 31
rect 7 28 9 30
rect 11 28 24 30
rect 7 27 24 28
rect 28 30 35 31
rect 28 28 30 30
rect 32 28 35 30
rect 28 27 35 28
rect 46 46 50 48
rect 46 44 47 46
rect 49 44 50 46
rect 46 30 50 44
rect 53 37 57 58
rect 69 58 75 60
rect 69 56 72 58
rect 74 56 75 58
rect 69 54 75 56
rect 69 47 73 54
rect 60 46 73 47
rect 60 44 62 46
rect 64 44 73 46
rect 120 61 126 69
rect 161 63 165 69
rect 182 67 184 69
rect 186 67 188 69
rect 182 66 188 67
rect 94 58 99 60
rect 120 59 122 61
rect 124 59 126 61
rect 120 58 126 59
rect 150 61 157 62
rect 150 59 152 61
rect 154 59 157 61
rect 161 61 162 63
rect 164 61 165 63
rect 161 59 165 61
rect 150 58 157 59
rect 94 56 95 58
rect 97 56 99 58
rect 94 54 99 56
rect 60 43 73 44
rect 53 35 54 37
rect 56 35 57 37
rect 53 33 57 35
rect 69 39 73 43
rect 69 37 75 39
rect 69 35 72 37
rect 74 35 75 37
rect 69 33 75 35
rect 95 30 99 54
rect 110 56 114 58
rect 110 54 111 56
rect 113 55 114 56
rect 131 56 135 58
rect 113 54 128 55
rect 110 51 128 54
rect 124 46 128 51
rect 124 44 125 46
rect 127 44 128 46
rect 124 39 128 44
rect 120 35 128 39
rect 131 54 132 56
rect 134 54 135 56
rect 120 31 124 35
rect 131 31 135 54
rect 46 29 99 30
rect 46 27 95 29
rect 97 27 99 29
rect 111 27 124 31
rect 128 30 135 31
rect 128 28 130 30
rect 132 28 135 30
rect 128 27 135 28
rect 46 26 99 27
rect 146 46 150 48
rect 146 44 147 46
rect 149 44 150 46
rect 146 30 150 44
rect 153 37 157 58
rect 169 58 175 60
rect 169 56 172 58
rect 174 56 175 58
rect 169 54 175 56
rect 169 47 173 54
rect 160 46 173 47
rect 160 44 162 46
rect 164 44 173 46
rect 220 61 226 69
rect 261 63 265 69
rect 282 67 284 69
rect 286 67 288 69
rect 282 66 288 67
rect 194 58 199 60
rect 220 59 222 61
rect 224 59 226 61
rect 220 58 226 59
rect 250 61 257 62
rect 250 59 252 61
rect 254 59 257 61
rect 261 61 262 63
rect 264 61 265 63
rect 261 59 265 61
rect 250 58 257 59
rect 194 56 195 58
rect 197 56 199 58
rect 194 54 199 56
rect 160 43 173 44
rect 153 35 154 37
rect 156 35 157 37
rect 153 33 157 35
rect 169 39 173 43
rect 169 37 175 39
rect 169 35 172 37
rect 174 35 175 37
rect 169 33 175 35
rect 195 30 199 54
rect 210 56 214 58
rect 210 54 211 56
rect 213 55 214 56
rect 231 56 235 58
rect 213 54 228 55
rect 210 51 228 54
rect 224 46 228 51
rect 224 44 225 46
rect 227 44 228 46
rect 224 39 228 44
rect 220 35 228 39
rect 231 54 232 56
rect 234 54 235 56
rect 220 31 224 35
rect 231 31 235 54
rect 146 29 199 30
rect 146 27 195 29
rect 197 27 199 29
rect 207 30 224 31
rect 207 28 209 30
rect 211 28 224 30
rect 207 27 224 28
rect 228 30 235 31
rect 228 28 230 30
rect 232 28 235 30
rect 228 27 235 28
rect 146 26 199 27
rect 246 46 250 48
rect 246 44 247 46
rect 249 44 250 46
rect 246 30 250 44
rect 253 37 257 58
rect 269 58 275 60
rect 269 56 272 58
rect 274 56 275 58
rect 269 54 275 56
rect 269 47 273 54
rect 260 46 273 47
rect 260 44 262 46
rect 264 44 273 46
rect 320 61 326 69
rect 361 63 365 69
rect 382 67 384 69
rect 386 67 388 69
rect 382 66 388 67
rect 294 58 299 60
rect 320 59 322 61
rect 324 59 326 61
rect 320 58 326 59
rect 350 61 357 62
rect 350 59 352 61
rect 354 59 357 61
rect 361 61 362 63
rect 364 61 365 63
rect 361 59 365 61
rect 350 58 357 59
rect 294 56 295 58
rect 297 56 299 58
rect 294 54 299 56
rect 260 43 273 44
rect 253 35 254 37
rect 256 35 257 37
rect 253 33 257 35
rect 269 39 273 43
rect 269 37 275 39
rect 269 35 272 37
rect 274 35 275 37
rect 269 33 275 35
rect 295 30 299 54
rect 310 56 314 58
rect 310 54 311 56
rect 313 55 314 56
rect 331 56 335 58
rect 313 54 328 55
rect 310 51 328 54
rect 324 46 328 51
rect 324 44 325 46
rect 327 44 328 46
rect 324 39 328 44
rect 320 35 328 39
rect 331 54 332 56
rect 334 54 335 56
rect 320 31 324 35
rect 331 31 335 54
rect 246 29 299 30
rect 246 27 295 29
rect 297 27 299 29
rect 307 30 324 31
rect 307 28 309 30
rect 311 28 324 30
rect 307 27 324 28
rect 328 30 335 31
rect 328 28 330 30
rect 332 28 335 30
rect 328 27 335 28
rect 246 26 299 27
rect 346 46 350 48
rect 346 44 347 46
rect 349 44 350 46
rect 346 30 350 44
rect 353 37 357 58
rect 369 58 375 60
rect 420 61 426 69
rect 461 63 465 69
rect 482 67 484 69
rect 486 67 488 69
rect 482 66 488 67
rect 369 56 372 58
rect 374 56 375 58
rect 369 54 375 56
rect 369 47 373 54
rect 394 58 399 60
rect 420 59 422 61
rect 424 59 426 61
rect 420 58 426 59
rect 450 61 457 62
rect 450 59 452 61
rect 454 59 457 61
rect 461 61 462 63
rect 464 61 465 63
rect 461 59 465 61
rect 450 58 457 59
rect 394 56 395 58
rect 397 56 399 58
rect 394 54 399 56
rect 360 46 373 47
rect 360 44 362 46
rect 364 44 373 46
rect 360 43 373 44
rect 353 35 354 37
rect 356 35 357 37
rect 353 33 357 35
rect 369 39 373 43
rect 369 37 375 39
rect 369 35 372 37
rect 374 35 375 37
rect 369 33 375 35
rect 395 30 399 54
rect 410 56 414 58
rect 410 54 411 56
rect 413 55 414 56
rect 431 56 435 58
rect 413 54 428 55
rect 410 51 428 54
rect 424 46 428 51
rect 424 44 425 46
rect 427 44 428 46
rect 424 39 428 44
rect 420 35 428 39
rect 431 54 432 56
rect 434 54 435 56
rect 420 31 424 35
rect 431 31 435 54
rect 346 29 399 30
rect 346 27 395 29
rect 397 27 399 29
rect 407 30 424 31
rect 407 28 409 30
rect 411 28 424 30
rect 407 27 424 28
rect 428 30 435 31
rect 428 28 430 30
rect 432 28 435 30
rect 428 27 435 28
rect 346 26 399 27
rect 446 46 450 48
rect 446 44 447 46
rect 449 44 450 46
rect 446 30 450 44
rect 453 37 457 58
rect 469 58 475 60
rect 469 56 472 58
rect 474 56 475 58
rect 469 54 475 56
rect 469 47 473 54
rect 494 58 499 60
rect 494 56 495 58
rect 497 56 499 58
rect 494 54 499 56
rect 460 46 473 47
rect 460 44 462 46
rect 464 44 473 46
rect 460 43 473 44
rect 453 35 454 37
rect 456 35 457 37
rect 453 33 457 35
rect 469 39 473 43
rect 469 37 475 39
rect 469 35 472 37
rect 474 35 475 37
rect 469 33 475 35
rect 495 30 499 54
rect 520 61 526 69
rect 561 63 565 69
rect 582 67 584 69
rect 586 67 588 69
rect 582 66 588 67
rect 520 59 522 61
rect 524 59 526 61
rect 520 58 526 59
rect 550 61 557 62
rect 550 59 552 61
rect 554 59 557 61
rect 561 61 562 63
rect 564 61 565 63
rect 561 59 565 61
rect 550 58 557 59
rect 510 56 514 58
rect 510 54 511 56
rect 513 55 514 56
rect 531 56 535 58
rect 513 54 528 55
rect 510 51 528 54
rect 524 46 528 51
rect 524 44 525 46
rect 527 44 528 46
rect 524 39 528 44
rect 520 35 528 39
rect 531 54 532 56
rect 534 54 535 56
rect 520 31 524 35
rect 531 31 535 54
rect 446 29 499 30
rect 446 27 495 29
rect 497 27 499 29
rect 507 30 524 31
rect 507 28 509 30
rect 511 28 524 30
rect 507 27 524 28
rect 528 30 535 31
rect 528 28 530 30
rect 532 28 535 30
rect 528 27 535 28
rect 446 26 499 27
rect 546 46 550 48
rect 546 44 547 46
rect 549 44 550 46
rect 546 30 550 44
rect 553 37 557 58
rect 569 58 575 60
rect 569 56 572 58
rect 574 56 575 58
rect 569 54 575 56
rect 569 47 573 54
rect 594 58 599 60
rect 594 56 595 58
rect 597 56 599 58
rect 594 54 599 56
rect 560 46 573 47
rect 560 44 562 46
rect 564 44 573 46
rect 560 43 573 44
rect 553 35 554 37
rect 556 35 557 37
rect 553 33 557 35
rect 569 39 573 43
rect 569 37 575 39
rect 569 35 572 37
rect 574 35 575 37
rect 569 33 575 35
rect 595 30 599 54
rect 620 61 626 69
rect 661 63 665 69
rect 682 67 684 69
rect 686 67 688 69
rect 682 66 688 67
rect 620 59 622 61
rect 624 59 626 61
rect 620 58 626 59
rect 650 61 657 62
rect 650 59 652 61
rect 654 59 657 61
rect 661 61 662 63
rect 664 61 665 63
rect 661 59 665 61
rect 650 58 657 59
rect 610 56 614 58
rect 610 54 611 56
rect 613 55 614 56
rect 631 56 635 58
rect 613 54 628 55
rect 610 51 628 54
rect 624 46 628 51
rect 624 44 625 46
rect 627 44 628 46
rect 624 39 628 44
rect 620 35 628 39
rect 631 54 632 56
rect 634 54 635 56
rect 620 31 624 35
rect 631 31 635 54
rect 546 29 599 30
rect 546 27 595 29
rect 597 27 599 29
rect 607 30 624 31
rect 607 28 609 30
rect 611 28 624 30
rect 607 27 624 28
rect 628 30 635 31
rect 628 28 630 30
rect 632 28 635 30
rect 628 27 635 28
rect 546 26 599 27
rect 646 46 650 48
rect 646 44 647 46
rect 649 44 650 46
rect 646 30 650 44
rect 653 37 657 58
rect 669 58 675 60
rect 669 56 672 58
rect 674 56 675 58
rect 669 54 675 56
rect 669 47 673 54
rect 694 58 699 60
rect 694 56 695 58
rect 697 56 699 58
rect 694 54 699 56
rect 660 46 673 47
rect 660 44 662 46
rect 664 44 673 46
rect 660 43 673 44
rect 653 35 654 37
rect 656 35 657 37
rect 653 33 657 35
rect 669 39 673 43
rect 669 37 675 39
rect 669 35 672 37
rect 674 35 675 37
rect 669 33 675 35
rect 695 30 699 54
rect 720 61 726 69
rect 761 63 765 69
rect 782 67 784 69
rect 786 67 788 69
rect 782 66 788 67
rect 720 59 722 61
rect 724 59 726 61
rect 720 58 726 59
rect 750 61 757 62
rect 750 59 752 61
rect 754 59 757 61
rect 761 61 762 63
rect 764 61 765 63
rect 761 59 765 61
rect 750 58 757 59
rect 710 56 714 58
rect 710 54 711 56
rect 713 55 714 56
rect 731 56 735 58
rect 713 54 728 55
rect 710 51 728 54
rect 724 46 728 51
rect 724 44 725 46
rect 727 44 728 46
rect 724 39 728 44
rect 720 35 728 39
rect 731 54 732 56
rect 734 54 735 56
rect 720 31 724 35
rect 731 31 735 54
rect 646 29 699 30
rect 646 27 695 29
rect 697 27 699 29
rect 707 30 724 31
rect 707 28 709 30
rect 711 28 724 30
rect 707 27 724 28
rect 728 30 735 31
rect 728 28 730 30
rect 732 28 735 30
rect 728 27 735 28
rect 646 26 699 27
rect 746 46 750 48
rect 746 44 747 46
rect 749 44 750 46
rect 746 30 750 44
rect 753 37 757 58
rect 769 58 775 60
rect 769 56 772 58
rect 774 56 775 58
rect 769 54 775 56
rect 769 47 773 54
rect 794 58 799 60
rect 794 56 795 58
rect 797 56 799 58
rect 794 54 799 56
rect 760 46 773 47
rect 760 44 762 46
rect 764 44 773 46
rect 760 43 773 44
rect 753 35 754 37
rect 756 35 757 37
rect 753 33 757 35
rect 769 39 773 43
rect 769 37 775 39
rect 769 35 772 37
rect 774 35 775 37
rect 769 33 775 35
rect 795 30 799 54
rect 746 29 799 30
rect 746 27 795 29
rect 797 27 799 29
rect 746 26 799 27
rect 18 22 24 23
rect 18 20 20 22
rect 22 20 24 22
rect 18 13 24 20
rect 118 22 124 23
rect 62 21 68 22
rect 62 19 64 21
rect 66 19 68 21
rect 62 13 68 19
rect 81 21 87 22
rect 81 19 83 21
rect 85 19 87 21
rect 81 13 87 19
rect 118 20 120 22
rect 122 20 124 22
rect 118 13 124 20
rect 218 22 224 23
rect 162 21 168 22
rect 162 19 164 21
rect 166 19 168 21
rect 162 13 168 19
rect 181 21 187 22
rect 181 19 183 21
rect 185 19 187 21
rect 181 13 187 19
rect 218 20 220 22
rect 222 20 224 22
rect 218 13 224 20
rect 318 22 324 23
rect 262 21 268 22
rect 262 19 264 21
rect 266 19 268 21
rect 262 13 268 19
rect 281 21 287 22
rect 281 19 283 21
rect 285 19 287 21
rect 281 13 287 19
rect 318 20 320 22
rect 322 20 324 22
rect 318 13 324 20
rect 418 22 424 23
rect 362 21 368 22
rect 362 19 364 21
rect 366 19 368 21
rect 362 13 368 19
rect 381 21 387 22
rect 381 19 383 21
rect 385 19 387 21
rect 381 13 387 19
rect 418 20 420 22
rect 422 20 424 22
rect 418 13 424 20
rect 518 22 524 23
rect 462 21 468 22
rect 462 19 464 21
rect 466 19 468 21
rect 462 13 468 19
rect 481 21 487 22
rect 481 19 483 21
rect 485 19 487 21
rect 481 13 487 19
rect 518 20 520 22
rect 522 20 524 22
rect 518 13 524 20
rect 618 22 624 23
rect 562 21 568 22
rect 562 19 564 21
rect 566 19 568 21
rect 562 13 568 19
rect 581 21 587 22
rect 581 19 583 21
rect 585 19 587 21
rect 581 13 587 19
rect 618 20 620 22
rect 622 20 624 22
rect 618 13 624 20
rect 718 22 724 23
rect 662 21 668 22
rect 662 19 664 21
rect 666 19 668 21
rect 662 13 668 19
rect 681 21 687 22
rect 681 19 683 21
rect 685 19 687 21
rect 681 13 687 19
rect 718 20 720 22
rect 722 20 724 22
rect 718 13 724 20
rect 762 21 768 22
rect 762 19 764 21
rect 766 19 768 21
rect 762 13 768 19
rect 781 21 787 22
rect 781 19 783 21
rect 785 19 787 21
rect 781 13 787 19
<< via1 >>
rect 8 323 10 325
rect 80 340 82 342
rect 180 348 182 350
rect 88 339 90 341
rect 108 324 110 326
rect 140 320 142 322
rect 188 339 190 341
rect 208 323 210 325
rect 240 327 242 329
rect 280 347 282 349
rect 288 339 290 341
rect 308 331 310 333
rect 340 323 342 325
rect 388 339 390 341
rect 388 323 390 325
rect 408 323 410 325
rect 440 319 442 321
rect 488 339 490 341
rect 480 329 482 331
rect 503 347 505 349
rect 540 331 542 333
rect 603 348 605 350
rect 588 339 590 341
rect 588 323 590 325
rect 640 331 642 333
rect 688 339 690 341
rect 688 323 690 325
rect 704 347 706 349
rect 788 339 790 341
rect 788 323 790 325
rect 31 308 33 310
rect 731 308 733 310
rect 24 254 26 256
rect 16 245 18 247
rect 65 237 67 239
rect 101 237 103 239
rect 116 262 118 264
rect 116 245 118 247
rect 201 261 203 263
rect 193 254 195 256
rect 224 254 226 256
rect 216 245 218 247
rect 165 237 167 239
rect 301 262 303 264
rect 316 262 318 264
rect 316 245 318 247
rect 265 237 267 239
rect 393 254 395 256
rect 365 237 367 239
rect 403 237 405 239
rect 426 254 428 256
rect 418 245 420 247
rect 503 262 505 264
rect 518 262 520 264
rect 518 245 520 247
rect 467 237 469 239
rect 595 254 597 256
rect 626 254 628 256
rect 618 245 620 247
rect 567 237 569 239
rect 703 262 705 264
rect 718 262 720 264
rect 718 245 720 247
rect 667 237 669 239
rect 795 254 797 256
rect 767 237 769 239
rect 16 195 18 197
rect 101 203 103 205
rect 16 179 18 181
rect 116 195 118 197
rect 124 187 126 189
rect 64 169 66 171
rect 196 179 198 181
rect 216 195 218 197
rect 300 204 302 206
rect 216 179 218 181
rect 296 187 298 189
rect 316 195 318 197
rect 324 187 326 189
rect 395 206 397 208
rect 395 179 397 181
rect 418 195 420 197
rect 418 179 420 181
rect 498 187 500 189
rect 518 195 520 197
rect 526 187 528 189
rect 598 179 600 181
rect 618 195 620 197
rect 618 179 620 181
rect 698 187 700 189
rect 718 195 720 197
rect 726 187 728 189
rect 813 189 815 191
rect 797 179 799 181
rect 173 164 175 166
rect 273 164 275 166
rect 373 164 375 166
rect 475 164 477 166
rect 575 164 577 166
rect 675 164 677 166
rect 775 164 777 166
rect 16 117 18 119
rect 64 113 66 115
rect 96 117 98 119
rect 124 109 126 111
rect 25 92 27 94
rect 264 128 266 130
rect 164 101 166 103
rect 200 117 202 119
rect 124 92 126 94
rect 224 101 226 103
rect 296 117 298 119
rect 296 109 298 111
rect 316 117 318 119
rect 224 92 226 94
rect 364 109 366 111
rect 396 117 398 119
rect 418 117 420 119
rect 324 92 326 94
rect 566 128 568 130
rect 666 128 668 130
rect 466 121 468 123
rect 498 117 500 119
rect 526 110 528 112
rect 426 92 428 94
rect 602 101 604 103
rect 618 118 620 120
rect 527 92 529 94
rect 703 117 705 119
rect 695 110 697 112
rect 627 92 629 94
rect 726 104 728 106
rect 766 96 768 98
rect 797 117 799 119
rect 813 117 815 119
rect 727 92 729 94
rect 8 35 10 37
rect 80 52 82 54
rect 180 60 182 62
rect 88 51 90 53
rect 108 36 110 38
rect 188 51 190 53
rect 208 35 210 37
rect 280 59 282 61
rect 288 51 290 53
rect 308 43 310 45
rect 388 51 390 53
rect 388 35 390 37
rect 408 35 410 37
rect 488 51 490 53
rect 480 41 482 43
rect 503 59 505 61
rect 508 43 510 45
rect 603 60 605 62
rect 588 51 590 53
rect 588 35 590 37
rect 688 51 690 53
rect 688 35 690 37
rect 704 59 706 61
rect 788 51 790 53
rect 788 35 790 37
<< via2 >>
rect 821 339 823 341
rect 300 327 302 329
rect 599 331 601 333
rect 640 326 642 328
rect 31 302 33 304
rect 140 313 142 315
rect 440 323 442 325
rect 340 318 342 320
rect 731 302 733 304
rect 340 286 342 288
rect 703 286 705 288
rect 201 270 203 272
rect 301 270 303 272
rect 498 262 500 264
rect 703 270 705 272
rect 599 254 601 256
rect 789 254 791 256
rect 101 233 103 235
rect 265 220 267 222
rect 403 230 405 232
rect 503 226 505 228
rect 567 226 569 228
rect 667 218 669 220
rect 767 219 769 221
rect 403 206 405 208
rect 813 219 815 221
rect 403 187 405 189
rect 503 187 505 189
rect 702 187 704 189
rect 203 179 205 181
rect 603 179 605 181
rect 200 164 202 166
rect 300 164 302 166
rect 403 164 405 166
rect 96 154 98 156
rect 703 164 705 166
rect 575 154 577 156
rect 775 154 777 156
rect 200 138 202 140
rect 96 135 98 137
rect 264 121 266 123
rect 300 117 302 119
rect 498 138 500 140
rect 352 109 354 111
rect 506 130 508 132
rect 466 109 468 111
rect 606 130 608 132
rect 703 136 705 138
rect 666 120 668 122
rect 813 154 815 156
rect 64 100 66 102
rect 208 101 210 103
rect 8 86 10 88
rect 404 84 406 86
rect 606 84 608 86
rect 466 67 468 69
rect 821 51 823 53
rect 208 43 210 45
rect 304 43 306 45
rect 404 35 406 37
rect 666 35 668 37
rect 352 14 354 16
<< labels >>
rlabel alu1 17 245 17 245 1 s2
rlabel alu1 117 245 117 245 1 s2
rlabel alu1 217 245 217 245 1 s2
rlabel alu1 317 245 317 245 1 s2
rlabel alu1 17 197 17 197 1 s1
rlabel alu1 117 197 117 197 1 s1
rlabel alu1 217 197 217 197 1 s1
rlabel alu1 317 197 317 197 1 s1
rlabel alu1 317 101 317 101 1 s0
rlabel alu1 217 101 217 101 1 s0
rlabel alu1 117 101 117 101 1 s0
rlabel alu1 17 101 17 101 1 s0
rlabel alu1 17 261 17 261 1 a10
rlabel alu1 65 257 65 257 1 z0
rlabel alu1 97 257 97 257 1 a00
rlabel alu1 165 257 165 257 1 z4
rlabel alu1 197 257 197 257 1 a04
rlabel alu1 117 261 117 261 1 a14
rlabel alu1 217 261 217 261 1 a12
rlabel alu1 265 257 265 257 1 z2
rlabel alu1 297 257 297 257 1 a02
rlabel alu1 317 261 317 261 1 a16
rlabel alu1 365 257 365 257 1 z6
rlabel alu1 397 257 397 257 1 a06
rlabel alu1 17 181 17 181 1 b10
rlabel alu1 65 185 65 185 1 y0
rlabel alu1 97 187 97 187 1 b00
rlabel alu1 117 181 117 181 1 b12
rlabel alu1 165 185 165 185 1 y2
rlabel alu1 197 185 197 185 1 b02
rlabel alu1 217 181 217 181 1 b14
rlabel alu1 265 185 265 185 1 y4
rlabel alu1 297 185 297 185 1 b04
rlabel alu1 317 181 317 181 1 b16
rlabel alu1 365 185 365 185 1 y6
rlabel alu1 397 185 397 185 1 b06
rlabel alu1 455 225 455 225 4 vss
rlabel alu1 455 153 455 153 2 vdd
rlabel alu1 455 81 455 81 4 vss
rlabel alu1 419 245 419 245 1 s2
rlabel alu1 519 245 519 245 1 s2
rlabel alu1 619 245 619 245 1 s2
rlabel alu1 719 245 719 245 1 s2
rlabel alu1 419 197 419 197 1 s1
rlabel alu1 519 197 519 197 1 s1
rlabel alu1 619 197 619 197 1 s1
rlabel alu1 719 197 719 197 1 s1
rlabel alu1 719 101 719 101 1 s0
rlabel alu1 619 101 619 101 1 s0
rlabel alu1 519 101 519 101 1 s0
rlabel alu1 419 101 419 101 1 s0
rlabel alu1 467 257 467 257 1 z1
rlabel alu1 499 257 499 257 1 a01
rlabel alu1 567 257 567 257 1 z5
rlabel alu1 599 257 599 257 1 a05
rlabel alu1 619 261 619 261 1 a13
rlabel alu1 667 257 667 257 1 z3
rlabel alu1 699 257 699 257 1 a03
rlabel alu1 719 261 719 261 1 a17
rlabel alu1 767 257 767 257 1 z7
rlabel alu1 799 257 799 257 1 a07
rlabel alu1 519 261 519 261 1 a15
rlabel alu1 419 261 419 261 1 a11
rlabel alu1 799 185 799 185 1 b07
rlabel alu1 767 185 767 185 1 y7
rlabel alu1 719 181 719 181 1 b17
rlabel alu1 699 185 699 185 1 b05
rlabel alu1 667 185 667 185 1 y5
rlabel alu1 620 181 620 181 1 b15
rlabel alu1 599 185 599 185 1 b03
rlabel alu1 567 185 567 185 1 y3
rlabel alu1 519 181 519 181 1 b13
rlabel alu1 419 181 419 181 1 b11
rlabel alu1 467 185 467 185 1 y1
rlabel alu1 499 185 499 185 1 b01
rlabel alu1 17 117 17 117 1 c10
rlabel alu1 65 113 65 113 1 x0
rlabel alu1 97 113 97 113 1 c00
rlabel alu1 117 117 117 117 1 c12
rlabel alu1 165 113 165 113 1 x2
rlabel alu1 197 113 197 113 1 c02
rlabel alu1 217 117 217 117 1 c13
rlabel alu1 265 113 265 113 1 x3
rlabel alu1 297 113 297 113 1 c03
rlabel alu1 317 117 317 117 1 c11
rlabel alu1 365 113 365 113 1 x1
rlabel alu1 397 113 397 113 1 c01
rlabel alu1 419 117 419 117 1 c16
rlabel alu1 467 113 467 113 1 x6
rlabel alu1 499 113 499 113 1 c06
rlabel alu1 519 117 519 117 1 c14
rlabel alu1 567 113 567 113 1 x4
rlabel alu1 619 117 619 117 1 c15
rlabel alu1 667 113 667 113 1 x5
rlabel alu1 699 113 699 113 1 c05
rlabel alu1 719 117 719 117 1 c17
rlabel alu1 767 113 767 113 1 x7
rlabel alu1 799 113 799 113 1 c07
rlabel alu1 455 287 455 287 1 vdd
rlabel alu2 599 113 599 113 1 c04
rlabel alu1 353 297 353 297 8 vdd
rlabel alu1 353 9 353 9 8 vdd
rlabel alu1 353 73 353 73 8 vss
rlabel alu1 41 329 41 329 1 q0
rlabel alu1 89 325 89 325 1 p10
rlabel alu1 141 329 141 329 1 q1
rlabel alu1 189 325 189 325 1 p11
rlabel alu1 241 329 241 329 1 q2
rlabel alu1 289 325 289 325 1 p12
rlabel alu1 341 329 341 329 1 q3
rlabel alu1 381 327 381 327 1 p13
rlabel alu1 441 329 441 329 1 q4
rlabel alu1 489 325 489 325 1 p14
rlabel alu1 541 329 541 329 1 q5
rlabel alu1 582 326 582 326 1 p15
rlabel alu1 641 329 641 329 1 q6
rlabel alu1 689 327 689 327 1 p16
rlabel alu1 741 329 741 329 1 q7
rlabel alu1 781 329 781 329 1 p17
rlabel alu1 9 41 9 41 1 r00
rlabel alu1 89 37 89 37 1 r10
rlabel alu1 109 41 109 41 1 r01
rlabel alu1 189 37 189 37 1 r11
rlabel alu1 209 41 209 41 1 r02
rlabel alu1 289 37 289 37 1 r12
rlabel alu1 309 41 309 41 1 r03
rlabel alu1 381 39 381 39 1 r13
rlabel alu1 409 41 409 41 1 r04
rlabel alu1 489 37 489 37 1 r14
rlabel alu1 509 41 509 41 1 r05
rlabel alu1 582 38 582 38 1 r15
rlabel alu1 609 41 609 41 1 r06
rlabel alu1 689 39 689 39 1 r16
rlabel alu1 709 41 709 41 1 r07
rlabel alu1 781 41 781 41 1 r17
rlabel via1 89 340 89 340 1 left_right
rlabel via1 89 52 89 52 1 left_right
rlabel alu1 41 42 41 42 1 out0
rlabel alu1 141 41 141 41 1 out1
rlabel alu1 241 42 241 42 1 out2
rlabel alu1 341 41 341 41 1 out3
rlabel alu1 441 41 441 41 1 out4
rlabel alu1 541 41 541 41 1 out5
rlabel alu1 641 42 641 42 1 out6
rlabel alu1 741 41 741 41 1 out7
rlabel alu1 353 361 353 361 8 vss
rlabel alu2 403 279 403 279 1 LR
rlabel alu1 9 330 9 330 1 i0
rlabel alu1 109 329 109 329 1 i1
rlabel alu1 209 330 209 330 1 i2
rlabel alu1 309 329 309 329 1 i3
rlabel alu1 409 329 409 329 1 i4
rlabel alu1 509 330 509 330 1 i5
rlabel alu1 609 330 609 330 1 i6
rlabel alu1 709 329 709 329 1 i7
<< end >>
